
module osc (
	clkout,
	oscena);	

	output		clkout;
	input		oscena;
endmodule
