module char_rom (
    input [10:0] address,
    input clock,
    output [7:0] q
);

reg[7:0] q_reg;
reg[7:0] q_reg_2;

assign q = q_reg_2;

always @(posedge clock) begin
    case (address)
        // -- NUL: code x00
        0000: q_reg <= 8'b00000000; // 0
        0001: q_reg <= 8'b00000000; // 1
        0002: q_reg <= 8'b00000000; // 2
        0003: q_reg <= 8'b00000000; // 3
        0004: q_reg <= 8'b00000000; // 4
        0005: q_reg <= 8'b00000000; // 5
        0006: q_reg <= 8'b00000000; // 6
        0007: q_reg <= 8'b00000000; // 7
        0008: q_reg <= 8'b00000000; // 8
        0009: q_reg <= 8'b00000000; // 9
        0010: q_reg <= 8'b00000000; // a
        0011: q_reg <= 8'b00000000; // b
        0012: q_reg <= 8'b00000000; // c
        0013: q_reg <= 8'b00000000; // d
        0014: q_reg <= 8'b00000000; // e
        0015: q_reg <= 8'b00000000; // f
        // -- SOH: code x01
        0016: q_reg <= 8'b00000000; // 0
        0017: q_reg <= 8'b00000000; // 1
        0018: q_reg <= 8'b01111110; // 2  ******
        0019: q_reg <= 8'b10000001; // 3 *      *
        0020: q_reg <= 8'b10100101; // 4 * *  * *
        0021: q_reg <= 8'b10000001; // 5 *      *
        0022: q_reg <= 8'b10000001; // 6 *      *
        0023: q_reg <= 8'b10111101; // 7 * **** *
        0024: q_reg <= 8'b10011001; // 8 *  **  *
        0025: q_reg <= 8'b10000001; // 9 *      *
        0026: q_reg <= 8'b10000001; // a *      *
        0027: q_reg <= 8'b01111110; // b  ******
        0028: q_reg <= 8'b00000000; // c
        0029: q_reg <= 8'b00000000; // d
        0030: q_reg <= 8'b00000000; // e
        0031: q_reg <= 8'b00000000; // f
        // -- STX: code x02
        0032: q_reg <= 8'b00000000; // 0
        0033: q_reg <= 8'b00000000; // 1
        0034: q_reg <= 8'b01111110; // 2  ******
        0035: q_reg <= 8'b11111111; // 3 ********
        0036: q_reg <= 8'b11011011; // 4 ** ** **
        0037: q_reg <= 8'b11111111; // 5 ********
        0038: q_reg <= 8'b11111111; // 6 ********
        0039: q_reg <= 8'b11000011; // 7 **    **
        0040: q_reg <= 8'b11100111; // 8 ***  ***
        0041: q_reg <= 8'b11111111; // 9 ********
        0042: q_reg <= 8'b11111111; // a ********
        0043: q_reg <= 8'b01111110; // b  ******
        0044: q_reg <= 8'b00000000; // c
        0045: q_reg <= 8'b00000000; // d
        0046: q_reg <= 8'b00000000; // e
        0047: q_reg <= 8'b00000000; // f
        // -- ETX: code x03
        0048: q_reg <= 8'b00000000; // 0
        0049: q_reg <= 8'b00000000; // 1
        0050: q_reg <= 8'b00000000; // 2
        0051: q_reg <= 8'b00000000; // 3
        0052: q_reg <= 8'b01101100; // 4  ** **
        0053: q_reg <= 8'b11111110; // 5 *******
        0054: q_reg <= 8'b11111110; // 6 *******
        0055: q_reg <= 8'b11111110; // 7 *******
        0056: q_reg <= 8'b11111110; // 8 *******
        0057: q_reg <= 8'b01111100; // 9  *****
        0058: q_reg <= 8'b00111000; // a   ***
        0059: q_reg <= 8'b00010000; // b    *
        0060: q_reg <= 8'b00000000; // c
        0061: q_reg <= 8'b00000000; // d
        0062: q_reg <= 8'b00000000; // e
        0063: q_reg <= 8'b00000000; // f
        // -- EOT: code x04
        0064: q_reg <= 8'b00000000; // 0
        0065: q_reg <= 8'b00000000; // 1
        0066: q_reg <= 8'b00000000; // 2
        0067: q_reg <= 8'b00000000; // 3
        0068: q_reg <= 8'b00010000; // 4    *
        0069: q_reg <= 8'b00111000; // 5   ***
        0070: q_reg <= 8'b01111100; // 6  *****
        0071: q_reg <= 8'b11111110; // 7 *******
        0072: q_reg <= 8'b01111100; // 8  *****
        0073: q_reg <= 8'b00111000; // 9   ***
        0074: q_reg <= 8'b00010000; // a    *
        0075: q_reg <= 8'b00000000; // b
        0076: q_reg <= 8'b00000000; // c
        0077: q_reg <= 8'b00000000; // d
        0078: q_reg <= 8'b00000000; // e
        0079: q_reg <= 8'b00000000; // f
        // -- ENQ: code x05
        0080: q_reg <= 8'b00000000; // 0
        0081: q_reg <= 8'b00000000; // 1
        0082: q_reg <= 8'b00000000; // 2
        0083: q_reg <= 8'b00011000; // 3    **
        0084: q_reg <= 8'b00111100; // 4   ****
        0085: q_reg <= 8'b00111100; // 5   ****
        0086: q_reg <= 8'b11100111; // 6 ***  ***
        0087: q_reg <= 8'b11100111; // 7 ***  ***
        0088: q_reg <= 8'b11100111; // 8 ***  ***
        0089: q_reg <= 8'b00011000; // 9    **
        0090: q_reg <= 8'b00011000; // a    **
        0091: q_reg <= 8'b00111100; // b   ****
        0092: q_reg <= 8'b00000000; // c
        0093: q_reg <= 8'b00000000; // d
        0094: q_reg <= 8'b00000000; // e
        0095: q_reg <= 8'b00000000; // f
        // -- ACK: code x06
        0096: q_reg <= 8'b00000000; // 0
        0097: q_reg <= 8'b00000000; // 1
        0098: q_reg <= 8'b00000000; // 2
        0099: q_reg <= 8'b00011000; // 3    **
        0100: q_reg <= 8'b00111100; // 4   ****
        0101: q_reg <= 8'b01111110; // 5  ******
        0102: q_reg <= 8'b11111111; // 6 ********
        0103: q_reg <= 8'b11111111; // 7 ********
        0104: q_reg <= 8'b01111110; // 8  ******
        0105: q_reg <= 8'b00011000; // 9    **
        0106: q_reg <= 8'b00011000; // a    **
        0107: q_reg <= 8'b00111100; // b   ****
        0108: q_reg <= 8'b00000000; // c
        0109: q_reg <= 8'b00000000; // d
        0110: q_reg <= 8'b00000000; // e
        0111: q_reg <= 8'b00000000; // f
        // -- BEL: code x07
        0112: q_reg <= 8'b00000000; // 0
        0113: q_reg <= 8'b00000000; // 1
        0114: q_reg <= 8'b00000000; // 2
        0115: q_reg <= 8'b00000000; // 3
        0116: q_reg <= 8'b00000000; // 4
        0117: q_reg <= 8'b00000000; // 5
        0118: q_reg <= 8'b00011000; // 6    **
        0119: q_reg <= 8'b00111100; // 7   ****
        0120: q_reg <= 8'b00111100; // 8   ****
        0121: q_reg <= 8'b00011000; // 9    **
        0122: q_reg <= 8'b00000000; // a
        0123: q_reg <= 8'b00000000; // b
        0124: q_reg <= 8'b00000000; // c
        0125: q_reg <= 8'b00000000; // d
        0126: q_reg <= 8'b00000000; // e
        0127: q_reg <= 8'b00000000; // f
        // -- BS: code x08
        0128: q_reg <= 8'b11111111; // 0 ********
        0129: q_reg <= 8'b11111111; // 1 ********
        0130: q_reg <= 8'b11111111; // 2 ********
        0131: q_reg <= 8'b11111111; // 3 ********
        0132: q_reg <= 8'b11111111; // 4 ********
        0133: q_reg <= 8'b11111111; // 5 ********
        0134: q_reg <= 8'b11100111; // 6 ***  ***
        0135: q_reg <= 8'b11000011; // 7 **    **
        0136: q_reg <= 8'b11000011; // 8 **    **
        0137: q_reg <= 8'b11100111; // 9 ***  ***
        0138: q_reg <= 8'b11111111; // a ********
        0139: q_reg <= 8'b11111111; // b ********
        0140: q_reg <= 8'b11111111; // c ********
        0141: q_reg <= 8'b11111111; // d ********
        0142: q_reg <= 8'b11111111; // e ********
        0143: q_reg <= 8'b11111111; // f ********
        // -- HT: code x09
        0144: q_reg <= 8'b00000000; // 0
        0145: q_reg <= 8'b00000000; // 1
        0146: q_reg <= 8'b00000000; // 2
        0147: q_reg <= 8'b00000000; // 3
        0148: q_reg <= 8'b00000000; // 4
        0149: q_reg <= 8'b00111100; // 5   ****
        0150: q_reg <= 8'b01100110; // 6  **  **
        0151: q_reg <= 8'b01000010; // 7  *    *
        0152: q_reg <= 8'b01000010; // 8  *    *
        0153: q_reg <= 8'b01100110; // 9  **  **
        0154: q_reg <= 8'b00111100; // a   ****
        0155: q_reg <= 8'b00000000; // b
        0156: q_reg <= 8'b00000000; // c
        0157: q_reg <= 8'b00000000; // d
        0158: q_reg <= 8'b00000000; // e
        0159: q_reg <= 8'b00000000; // f
        // -- LF: code x0a
        0160: q_reg <= 8'b11111111; // 0 ********
        0161: q_reg <= 8'b11111111; // 1 ********
        0162: q_reg <= 8'b11111111; // 2 ********
        0163: q_reg <= 8'b11111111; // 3 ********
        0164: q_reg <= 8'b11111111; // 4 ********
        0165: q_reg <= 8'b11000011; // 5 **    **
        0166: q_reg <= 8'b10011001; // 6 *  **  *
        0167: q_reg <= 8'b10111101; // 7 * **** *
        0168: q_reg <= 8'b10111101; // 8 * **** *
        0169: q_reg <= 8'b10011001; // 9 *  **  *
        0170: q_reg <= 8'b11000011; // a **    **
        0171: q_reg <= 8'b11111111; // b ********
        0172: q_reg <= 8'b11111111; // c ********
        0173: q_reg <= 8'b11111111; // d ********
        0174: q_reg <= 8'b11111111; // e ********
        0175: q_reg <= 8'b11111111; // f ********
        // -- code x0b
        0176: q_reg <= 8'b00000000; // 0
        0177: q_reg <= 8'b00000000; // 1
        0178: q_reg <= 8'b00011110; // 2    ****
        0179: q_reg <= 8'b00001110; // 3     ***
        0180: q_reg <= 8'b00011010; // 4    ** *
        0181: q_reg <= 8'b00110010; // 5   **  *
        0182: q_reg <= 8'b01111000; // 6  ****
        0183: q_reg <= 8'b11001100; // 7 **  **
        0184: q_reg <= 8'b11001100; // 8 **  **
        0185: q_reg <= 8'b11001100; // 9 **  **
        0186: q_reg <= 8'b11001100; // a **  **
        0187: q_reg <= 8'b01111000; // b  ****
        0188: q_reg <= 8'b00000000; // c
        0189: q_reg <= 8'b00000000; // d
        0190: q_reg <= 8'b00000000; // e
        0191: q_reg <= 8'b00000000; // f
        // -- code x0c
        0192: q_reg <= 8'b00000000; // 0
        0193: q_reg <= 8'b00000000; // 1
        0194: q_reg <= 8'b00111100; // 2   ****
        0195: q_reg <= 8'b01100110; // 3  **  **
        0196: q_reg <= 8'b01100110; // 4  **  **
        0197: q_reg <= 8'b01100110; // 5  **  **
        0198: q_reg <= 8'b01100110; // 6  **  **
        0199: q_reg <= 8'b00111100; // 7   ****
        0200: q_reg <= 8'b00011000; // 8    **
        0201: q_reg <= 8'b01111110; // 9  ******
        0202: q_reg <= 8'b00011000; // a    **
        0203: q_reg <= 8'b00011000; // b    **
        0204: q_reg <= 8'b00000000; // c
        0205: q_reg <= 8'b00000000; // d
        0206: q_reg <= 8'b00000000; // e
        0207: q_reg <= 8'b00000000; // f
        // -- code x0d
        0208: q_reg <= 8'b00000000; // 0
        0209: q_reg <= 8'b00000000; // 1
        0210: q_reg <= 8'b00111111; // 2   ******
        0211: q_reg <= 8'b00110011; // 3   **  **
        0212: q_reg <= 8'b00111111; // 4   ******
        0213: q_reg <= 8'b00110000; // 5   **
        0214: q_reg <= 8'b00110000; // 6   **
        0215: q_reg <= 8'b00110000; // 7   **
        0216: q_reg <= 8'b00110000; // 8   **
        0217: q_reg <= 8'b01110000; // 9  ***
        0218: q_reg <= 8'b11110000; // a ****
        0219: q_reg <= 8'b11100000; // b ***
        0220: q_reg <= 8'b00000000; // c
        0221: q_reg <= 8'b00000000; // d
        0222: q_reg <= 8'b00000000; // e
        0223: q_reg <= 8'b00000000; // f
        // -- code x0e
        0224: q_reg <= 8'b00000000; // 0
        0225: q_reg <= 8'b00000000; // 1
        0226: q_reg <= 8'b01111111; // 2  *******
        0227: q_reg <= 8'b01100011; // 3  **   **
        0228: q_reg <= 8'b01111111; // 4  *******
        0229: q_reg <= 8'b01100011; // 5  **   **
        0230: q_reg <= 8'b01100011; // 6  **   **
        0231: q_reg <= 8'b01100011; // 7  **   **
        0232: q_reg <= 8'b01100011; // 8  **   **
        0233: q_reg <= 8'b01100111; // 9  **  ***
        0234: q_reg <= 8'b11100111; // a ***  ***
        0235: q_reg <= 8'b11100110; // b ***  **
        0236: q_reg <= 8'b11000000; // c **
        0237: q_reg <= 8'b00000000; // d
        0238: q_reg <= 8'b00000000; // e
        0239: q_reg <= 8'b00000000; // f
        // -- code x0f
        0240: q_reg <= 8'b00000000; // 0
        0241: q_reg <= 8'b00000000; // 1
        0242: q_reg <= 8'b00000000; // 2
        0243: q_reg <= 8'b00011000; // 3    **
        0244: q_reg <= 8'b00011000; // 4    **
        0245: q_reg <= 8'b11011011; // 5 ** ** **
        0246: q_reg <= 8'b00111100; // 6   ****
        0247: q_reg <= 8'b11100111; // 7 ***  ***
        0248: q_reg <= 8'b00111100; // 8   ****
        0249: q_reg <= 8'b11011011; // 9 ** ** **
        0250: q_reg <= 8'b00011000; // a    **
        0251: q_reg <= 8'b00011000; // b    **
        0252: q_reg <= 8'b00000000; // c
        0253: q_reg <= 8'b00000000; // d
        0254: q_reg <= 8'b00000000; // e
        0255: q_reg <= 8'b00000000; // f
        // -- code x10
        0256: q_reg <= 8'b00000000; // 0
        0257: q_reg <= 8'b10000000; // 1 *
        0258: q_reg <= 8'b11000000; // 2 **
        0259: q_reg <= 8'b11100000; // 3 ***
        0260: q_reg <= 8'b11110000; // 4 ****
        0261: q_reg <= 8'b11111000; // 5 *****
        0262: q_reg <= 8'b11111110; // 6 *******
        0263: q_reg <= 8'b11111000; // 7 *****
        0264: q_reg <= 8'b11110000; // 8 ****
        0265: q_reg <= 8'b11100000; // 9 ***
        0266: q_reg <= 8'b11000000; // a **
        0267: q_reg <= 8'b10000000; // b *
        0268: q_reg <= 8'b00000000; // c
        0269: q_reg <= 8'b00000000; // d
        0270: q_reg <= 8'b00000000; // e
        0271: q_reg <= 8'b00000000; // f
        // -- code x11
        0272: q_reg <= 8'b00000000; // 0
        0273: q_reg <= 8'b00000010; // 1       *
        0274: q_reg <= 8'b00000110; // 2      **
        0275: q_reg <= 8'b00001110; // 3     ***
        0276: q_reg <= 8'b00011110; // 4    ****
        0277: q_reg <= 8'b00111110; // 5   *****
        0278: q_reg <= 8'b11111110; // 6 *******
        0279: q_reg <= 8'b00111110; // 7   *****
        0280: q_reg <= 8'b00011110; // 8    ****
        0281: q_reg <= 8'b00001110; // 9     ***
        0282: q_reg <= 8'b00000110; // a      **
        0283: q_reg <= 8'b00000010; // b       *
        0284: q_reg <= 8'b00000000; // c
        0285: q_reg <= 8'b00000000; // d
        0286: q_reg <= 8'b00000000; // e
        0287: q_reg <= 8'b00000000; // f
        // -- code x12
        0288: q_reg <= 8'b00000000; // 0
        0289: q_reg <= 8'b00000000; // 1
        0290: q_reg <= 8'b00011000; // 2    **
        0291: q_reg <= 8'b00111100; // 3   ****
        0292: q_reg <= 8'b01111110; // 4  ******
        0293: q_reg <= 8'b00011000; // 5    **
        0294: q_reg <= 8'b00011000; // 6    **
        0295: q_reg <= 8'b00011000; // 7    **
        0296: q_reg <= 8'b01111110; // 8  ******
        0297: q_reg <= 8'b00111100; // 9   ****
        0298: q_reg <= 8'b00011000; // a    **
        0299: q_reg <= 8'b00000000; // b
        0300: q_reg <= 8'b00000000; // c
        0301: q_reg <= 8'b00000000; // d
        0302: q_reg <= 8'b00000000; // e
        0303: q_reg <= 8'b00000000; // f
        // -- code x13 reassigned to special forward slash
        0304: q_reg <= 8'b00000001; // 0        *
        0305: q_reg <= 8'b00000001; // 1        *
        0306: q_reg <= 8'b00000010; // 2       *
        0307: q_reg <= 8'b00000010; // 3       *
        0308: q_reg <= 8'b00000100; // 4      *
        0309: q_reg <= 8'b00000100; // 5      *
        0310: q_reg <= 8'b00001000; // 6     *
        0311: q_reg <= 8'b00001000; // 7     *
        0312: q_reg <= 8'b00010000; // 8    *
        0313: q_reg <= 8'b00010000; // 9    *
        0314: q_reg <= 8'b00100000; // a   *
        0315: q_reg <= 8'b00100000; // b   *
        0316: q_reg <= 8'b01000000; // c  *
        0317: q_reg <= 8'b01000000; // d  *
        0318: q_reg <= 8'b10000000; // e *
        0319: q_reg <= 8'b10000000; // f *
        // -- code x14
        0320: q_reg <= 8'b00000000; // 0
        0321: q_reg <= 8'b00000000; // 1
        0322: q_reg <= 8'b00000000; // 2
        0323: q_reg <= 8'b00000000; // 3
        0324: q_reg <= 8'b00000000; // 4
        0325: q_reg <= 8'b00000000; // 5
        0326: q_reg <= 8'b00000000; // 6
        0327: q_reg <= 8'b00000000; // 7
        0328: q_reg <= 8'b00000000; // 8
        0329: q_reg <= 8'b00000000; // 9
        0330: q_reg <= 8'b00000000; // a
        0331: q_reg <= 8'b00000000; // b
        0332: q_reg <= 8'b00000000; // c
        0333: q_reg <= 8'b00000000; // d
        0334: q_reg <= 8'b00000000; // e
        0335: q_reg <= 8'b11111111; // f ********
        // -- code x15
        0336: q_reg <= 8'b10000000; // 0 *
        0337: q_reg <= 8'b10000000; // 1 *
        0338: q_reg <= 8'b01000000; // 2  *
        0339: q_reg <= 8'b01000000; // 3  *
        0340: q_reg <= 8'b00100000; // 4   *
        0341: q_reg <= 8'b00100000; // 5   *
        0342: q_reg <= 8'b00010000; // 6    *
        0343: q_reg <= 8'b00010000; // 7    *
        0344: q_reg <= 8'b00001000; // 8     *
        0345: q_reg <= 8'b00001000; // 9     *
        0346: q_reg <= 8'b00000100; // a      *
        0347: q_reg <= 8'b00000100; // b      *
        0348: q_reg <= 8'b00000010; // c       *
        0349: q_reg <= 8'b00000010; // d       *
        0350: q_reg <= 8'b00000001; // e        *
        0351: q_reg <= 8'b00000001; // f        *
        // -- code x16
        0352: q_reg <= 8'b00000001; // 0        *
        0353: q_reg <= 8'b00000001; // 1        *
        0354: q_reg <= 8'b00000010; // 2       *
        0355: q_reg <= 8'b00000010; // 3       *
        0356: q_reg <= 8'b00000100; // 4      *
        0357: q_reg <= 8'b00000100; // 5      *
        0358: q_reg <= 8'b00001000; // 6     *
        0359: q_reg <= 8'b00001000; // 7     *
        0360: q_reg <= 8'b00010000; // 8    *
        0361: q_reg <= 8'b00010000; // 9    *
        0362: q_reg <= 8'b00100000; // a   *
        0363: q_reg <= 8'b00100000; // b   *
        0364: q_reg <= 8'b01000000; // c  *
        0365: q_reg <= 8'b01000000; // d  *
        0366: q_reg <= 8'b10000000; // e *
        0367: q_reg <= 8'b11111111; // f ********
        // -- code x17
        0368: q_reg <= 8'b00000000; // 0 
        0369: q_reg <= 8'b10000000; // 1 *
        0370: q_reg <= 8'b01000000; // 2  *
        0371: q_reg <= 8'b00100000; // 3   *
        0372: q_reg <= 8'b00010011; // 4    *  **
        0373: q_reg <= 8'b00001100; // 5     **
        0374: q_reg <= 8'b00000000; // 6
        0375: q_reg <= 8'b00000000; // 7
        0376: q_reg <= 8'b00000000; // 8
        0377: q_reg <= 8'b00000000; // 9
        0378: q_reg <= 8'b00000000; // a
        0379: q_reg <= 8'b00000000; // b
        0380: q_reg <= 8'b00000000; // c
        0381: q_reg <= 8'b00000000; // d
        0382: q_reg <= 8'b00000000; // e
        0383: q_reg <= 8'b00000000; // f
        // -- code x18
        0384: q_reg <= 8'b00000011; // 0       **
        0385: q_reg <= 8'b00001101; // 1     ** *
        0386: q_reg <= 8'b00110010; // 2   **  *
        0387: q_reg <= 8'b11000010; // 3 **    *
        0388: q_reg <= 8'b00000100; // 4      *
        0389: q_reg <= 8'b00000100; // 5      *
        0390: q_reg <= 8'b00001000; // 6     *
        0391: q_reg <= 8'b00001000; // 7     *
        0392: q_reg <= 8'b00010000; // 8    *
        0393: q_reg <= 8'b00010000; // 9    *
        0394: q_reg <= 8'b00100000; // a   *
        0395: q_reg <= 8'b00100000; // b   *
        0396: q_reg <= 8'b01000000; // c  *
        0397: q_reg <= 8'b01000000; // d  *
        0398: q_reg <= 8'b10000000; // e *
        0399: q_reg <= 8'b10000000; // f *
        // -- code x19
        0400: q_reg <= 8'b00000000; // 0
        0401: q_reg <= 8'b00000000; // 1
        0402: q_reg <= 8'b00011000; // 2    **
        0403: q_reg <= 8'b00011000; // 3    **
        0404: q_reg <= 8'b00011000; // 4    **
        0405: q_reg <= 8'b00011000; // 5    **
        0406: q_reg <= 8'b00011000; // 6    **
        0407: q_reg <= 8'b00011000; // 7    **
        0408: q_reg <= 8'b00011000; // 8    **
        0409: q_reg <= 8'b01111110; // 9  ******
        0410: q_reg <= 8'b00111100; // a   ****
        0411: q_reg <= 8'b00011000; // b    **
        0412: q_reg <= 8'b00000000; // c
        0413: q_reg <= 8'b00000000; // d
        0414: q_reg <= 8'b00000000; // e
        0415: q_reg <= 8'b00000000; // f
        // -- code x1a
        0416: q_reg <= 8'b00000000; // 0
        0417: q_reg <= 8'b00000000; // 1
        0418: q_reg <= 8'b00000000; // 2
        0419: q_reg <= 8'b00000000; // 3
        0420: q_reg <= 8'b00000000; // 4
        0421: q_reg <= 8'b00011000; // 5    **
        0422: q_reg <= 8'b00001100; // 6     **
        0423: q_reg <= 8'b11111110; // 7 *******
        0424: q_reg <= 8'b00001100; // 8     **
        0425: q_reg <= 8'b00011000; // 9    **
        0426: q_reg <= 8'b00000000; // a
        0427: q_reg <= 8'b00000000; // b
        0428: q_reg <= 8'b00000000; // c
        0429: q_reg <= 8'b00000000; // d
        0430: q_reg <= 8'b00000000; // e
        0431: q_reg <= 8'b00000000; // f
        // -- code x1b
        0432: q_reg <= 8'b00000000; // 0
        0433: q_reg <= 8'b00000000; // 1
        0434: q_reg <= 8'b00000000; // 2
        0435: q_reg <= 8'b00000000; // 3
        0436: q_reg <= 8'b00000000; // 4
        0437: q_reg <= 8'b00110000; // 5   **
        0438: q_reg <= 8'b01100000; // 6  **
        0439: q_reg <= 8'b11111110; // 7 *******
        0440: q_reg <= 8'b01100000; // 8  **
        0441: q_reg <= 8'b00110000; // 9   **
        0442: q_reg <= 8'b00000000; // a
        0443: q_reg <= 8'b00000000; // b
        0444: q_reg <= 8'b00000000; // c
        0445: q_reg <= 8'b00000000; // d
        0446: q_reg <= 8'b00000000; // e
        0447: q_reg <= 8'b00000000; // f
        // -- code x1c
        0448: q_reg <= 8'b00000000; // 0
        0449: q_reg <= 8'b00000000; // 1
        0450: q_reg <= 8'b00000000; // 2
        0451: q_reg <= 8'b00000000; // 3
        0452: q_reg <= 8'b00000000; // 4
        0453: q_reg <= 8'b00000000; // 5
        0454: q_reg <= 8'b11000000; // 6 **
        0455: q_reg <= 8'b11000000; // 7 **
        0456: q_reg <= 8'b11000000; // 8 **
        0457: q_reg <= 8'b11111110; // 9 *******
        0458: q_reg <= 8'b00000000; // a
        0459: q_reg <= 8'b00000000; // b
        0460: q_reg <= 8'b00000000; // c
        0461: q_reg <= 8'b00000000; // d
        0462: q_reg <= 8'b00000000; // e
        0463: q_reg <= 8'b00000000; // f
        // -- code x1d
        0464: q_reg <= 8'b00000000; // 0
        0465: q_reg <= 8'b00000000; // 1
        0466: q_reg <= 8'b00000000; // 2
        0467: q_reg <= 8'b00000000; // 3
        0468: q_reg <= 8'b00000000; // 4
        0469: q_reg <= 8'b00100100; // 5   *  *
        0470: q_reg <= 8'b01100110; // 6  **  **
        0471: q_reg <= 8'b11111111; // 7 ********
        0472: q_reg <= 8'b01100110; // 8  **  **
        0473: q_reg <= 8'b00100100; // 9   *  *
        0474: q_reg <= 8'b00000000; // a
        0475: q_reg <= 8'b00000000; // b
        0476: q_reg <= 8'b00000000; // c
        0477: q_reg <= 8'b00000000; // d
        0478: q_reg <= 8'b00000000; // e
        0479: q_reg <= 8'b00000000; // f
        // -- code x1e
        0480: q_reg <= 8'b00000000; // 0
        0481: q_reg <= 8'b00000000; // 1
        0482: q_reg <= 8'b00000000; // 2
        0483: q_reg <= 8'b00000000; // 3
        0484: q_reg <= 8'b00010000; // 4    *
        0485: q_reg <= 8'b00111000; // 5   ***
        0486: q_reg <= 8'b00111000; // 6   ***
        0487: q_reg <= 8'b01111100; // 7  *****
        0488: q_reg <= 8'b01111100; // 8  *****
        0489: q_reg <= 8'b11111110; // 9 *******
        0490: q_reg <= 8'b11111110; // a *******
        0491: q_reg <= 8'b00000000; // b
        0492: q_reg <= 8'b00000000; // c
        0493: q_reg <= 8'b00000000; // d
        0494: q_reg <= 8'b00000000; // e
        0495: q_reg <= 8'b00000000; // f
        // -- code x1f
        0496: q_reg <= 8'b00000000; // 0
        0497: q_reg <= 8'b00000000; // 1
        0498: q_reg <= 8'b00000000; // 2
        0499: q_reg <= 8'b00000000; // 3
        0500: q_reg <= 8'b11111110; // 4 *******
        0501: q_reg <= 8'b11111110; // 5 *******
        0502: q_reg <= 8'b01111100; // 6  *****
        0503: q_reg <= 8'b01111100; // 7  *****
        0504: q_reg <= 8'b00111000; // 8   ***
        0505: q_reg <= 8'b00111000; // 9   ***
        0506: q_reg <= 8'b00010000; // a    *
        0507: q_reg <= 8'b00000000; // b
        0508: q_reg <= 8'b00000000; // c
        0509: q_reg <= 8'b00000000; // d
        0510: q_reg <= 8'b00000000; // e
        0511: q_reg <= 8'b00000000; // f
        // -- code x20
        0512: q_reg <= 8'b00000000; // 0
        0513: q_reg <= 8'b00000000; // 1
        0514: q_reg <= 8'b00000000; // 2
        0515: q_reg <= 8'b00000000; // 3
        0516: q_reg <= 8'b00000000; // 4
        0517: q_reg <= 8'b00000000; // 5
        0518: q_reg <= 8'b00000000; // 6
        0519: q_reg <= 8'b00000000; // 7
        0520: q_reg <= 8'b00000000; // 8
        0521: q_reg <= 8'b00000000; // 9
        0522: q_reg <= 8'b00000000; // a
        0523: q_reg <= 8'b00000000; // b
        0524: q_reg <= 8'b00000000; // c
        0525: q_reg <= 8'b00000000; // d
        0526: q_reg <= 8'b00000000; // e
        0527: q_reg <= 8'b00000000; // f
        // -- code x21
        0528: q_reg <= 8'b00000000; // 0
        0529: q_reg <= 8'b00000000; // 1
        0530: q_reg <= 8'b00011000; // 2    **
        0531: q_reg <= 8'b00111100; // 3   ****
        0532: q_reg <= 8'b00111100; // 4   ****
        0533: q_reg <= 8'b00111100; // 5   ****
        0534: q_reg <= 8'b00011000; // 6    **
        0535: q_reg <= 8'b00011000; // 7    **
        0536: q_reg <= 8'b00011000; // 8    **
        0537: q_reg <= 8'b00000000; // 9
        0538: q_reg <= 8'b00011000; // a    **
        0539: q_reg <= 8'b00011000; // b    **
        0540: q_reg <= 8'b00000000; // c
        0541: q_reg <= 8'b00000000; // d
        0542: q_reg <= 8'b00000000; // e
        0543: q_reg <= 8'b00000000; // f
        // -- code x22
        0544: q_reg <= 8'b00000000; // 0
        0545: q_reg <= 8'b01100110; // 1  **  **
        0546: q_reg <= 8'b01100110; // 2  **  **
        0547: q_reg <= 8'b01100110; // 3  **  **
        0548: q_reg <= 8'b00100100; // 4   *  *
        0549: q_reg <= 8'b00000000; // 5
        0550: q_reg <= 8'b00000000; // 6
        0551: q_reg <= 8'b00000000; // 7
        0552: q_reg <= 8'b00000000; // 8
        0553: q_reg <= 8'b00000000; // 9
        0554: q_reg <= 8'b00000000; // a
        0555: q_reg <= 8'b00000000; // b
        0556: q_reg <= 8'b00000000; // c
        0557: q_reg <= 8'b00000000; // d
        0558: q_reg <= 8'b00000000; // e
        0559: q_reg <= 8'b00000000; // f
        // -- code x23
        0560: q_reg <= 8'b00000000; // 0
        0561: q_reg <= 8'b00000000; // 1
        0562: q_reg <= 8'b00000000; // 2
        0563: q_reg <= 8'b01101100; // 3  ** **
        0564: q_reg <= 8'b01101100; // 4  ** **
        0565: q_reg <= 8'b11111110; // 5 *******
        0566: q_reg <= 8'b01101100; // 6  ** **
        0567: q_reg <= 8'b01101100; // 7  ** **
        0568: q_reg <= 8'b01101100; // 8  ** **
        0569: q_reg <= 8'b11111110; // 9 *******
        0570: q_reg <= 8'b01101100; // a  ** **
        0571: q_reg <= 8'b01101100; // b  ** **
        0572: q_reg <= 8'b00000000; // c
        0573: q_reg <= 8'b00000000; // d
        0574: q_reg <= 8'b00000000; // e
        0575: q_reg <= 8'b00000000; // f
        // -- code x24
        0576: q_reg <= 8'b00011000; // 0     **
        0577: q_reg <= 8'b00011000; // 1     **
        0578: q_reg <= 8'b01111100; // 2   *****
        0579: q_reg <= 8'b11000110; // 3  **   **
        0580: q_reg <= 8'b11000010; // 4  **    *
        0581: q_reg <= 8'b11000000; // 5  **
        0582: q_reg <= 8'b01111100; // 6   *****
        0583: q_reg <= 8'b00000110; // 7       **
        0584: q_reg <= 8'b00000110; // 8       **
        0585: q_reg <= 8'b10000110; // 9  *    **
        0586: q_reg <= 8'b11000110; // a  **   **
        0587: q_reg <= 8'b01111100; // b   *****
        0588: q_reg <= 8'b00011000; // c     **
        0589: q_reg <= 8'b00011000; // d     **
        0590: q_reg <= 8'b00000000; // e
        0591: q_reg <= 8'b00000000; // f
        // -- code x25
        0592: q_reg <= 8'b00000000; // 0
        0593: q_reg <= 8'b00000000; // 1
        0594: q_reg <= 8'b00000000; // 2
        0595: q_reg <= 8'b00000000; // 3
        0596: q_reg <= 8'b11000010; // 4 **    *
        0597: q_reg <= 8'b11000110; // 5 **   **
        0598: q_reg <= 8'b00001100; // 6     **
        0599: q_reg <= 8'b00011000; // 7    **
        0600: q_reg <= 8'b00110000; // 8   **
        0601: q_reg <= 8'b01100000; // 9  **
        0602: q_reg <= 8'b11000110; // a **   **
        0603: q_reg <= 8'b10000110; // b *    **
        0604: q_reg <= 8'b00000000; // c
        0605: q_reg <= 8'b00000000; // d
        0606: q_reg <= 8'b00000000; // e
        0607: q_reg <= 8'b00000000; // f
        // -- code x26
        0608: q_reg <= 8'b00000000; // 0
        0609: q_reg <= 8'b00000000; // 1
        0610: q_reg <= 8'b00111000; // 2   ***
        0611: q_reg <= 8'b01101100; // 3  ** **
        0612: q_reg <= 8'b01101100; // 4  ** **
        0613: q_reg <= 8'b00111000; // 5   ***
        0614: q_reg <= 8'b01110110; // 6  *** **
        0615: q_reg <= 8'b11011100; // 7 ** ***
        0616: q_reg <= 8'b11001100; // 8 **  **
        0617: q_reg <= 8'b11001100; // 9 **  **
        0618: q_reg <= 8'b11001100; // a **  **
        0619: q_reg <= 8'b01110110; // b  *** **
        0620: q_reg <= 8'b00000000; // c
        0621: q_reg <= 8'b00000000; // d
        0622: q_reg <= 8'b00000000; // e
        0623: q_reg <= 8'b00000000; // f
        // -- code x27
        0624: q_reg <= 8'b00000000; // 0
        0625: q_reg <= 8'b00110000; // 1   **
        0626: q_reg <= 8'b00110000; // 2   **
        0627: q_reg <= 8'b00110000; // 3   **
        0628: q_reg <= 8'b01100000; // 4  **
        0629: q_reg <= 8'b00000000; // 5
        0630: q_reg <= 8'b00000000; // 6
        0631: q_reg <= 8'b00000000; // 7
        0632: q_reg <= 8'b00000000; // 8
        0633: q_reg <= 8'b00000000; // 9
        0634: q_reg <= 8'b00000000; // a
        0635: q_reg <= 8'b00000000; // b
        0636: q_reg <= 8'b00000000; // c
        0637: q_reg <= 8'b00000000; // d
        0638: q_reg <= 8'b00000000; // e
        0639: q_reg <= 8'b00000000; // f
        // -- code x28
        0640: q_reg <= 8'b00000000; // 0
        0641: q_reg <= 8'b00000000; // 1
        0642: q_reg <= 8'b00001100; // 2     **
        0643: q_reg <= 8'b00011000; // 3    **
        0644: q_reg <= 8'b00110000; // 4   **
        0645: q_reg <= 8'b00110000; // 5   **
        0646: q_reg <= 8'b00110000; // 6   **
        0647: q_reg <= 8'b00110000; // 7   **
        0648: q_reg <= 8'b00110000; // 8   **
        0649: q_reg <= 8'b00110000; // 9   **
        0650: q_reg <= 8'b00011000; // a    **
        0651: q_reg <= 8'b00001100; // b     **
        0652: q_reg <= 8'b00000000; // c
        0653: q_reg <= 8'b00000000; // d
        0654: q_reg <= 8'b00000000; // e
        0655: q_reg <= 8'b00000000; // f
        // -- code x29
        0656: q_reg <= 8'b00000000; // 0
        0657: q_reg <= 8'b00000000; // 1
        0658: q_reg <= 8'b00110000; // 2   **
        0659: q_reg <= 8'b00011000; // 3    **
        0660: q_reg <= 8'b00001100; // 4     **
        0661: q_reg <= 8'b00001100; // 5     **
        0662: q_reg <= 8'b00001100; // 6     **
        0663: q_reg <= 8'b00001100; // 7     **
        0664: q_reg <= 8'b00001100; // 8     **
        0665: q_reg <= 8'b00001100; // 9     **
        0666: q_reg <= 8'b00011000; // a    **
        0667: q_reg <= 8'b00110000; // b   **
        0668: q_reg <= 8'b00000000; // c
        0669: q_reg <= 8'b00000000; // d
        0670: q_reg <= 8'b00000000; // e
        0671: q_reg <= 8'b00000000; // f
        // -- code x2a
        0672: q_reg <= 8'b00000000; // 0
        0673: q_reg <= 8'b00000000; // 1
        0674: q_reg <= 8'b00000000; // 2
        0675: q_reg <= 8'b00000000; // 3
        0676: q_reg <= 8'b00000000; // 4
        0677: q_reg <= 8'b01100110; // 5  **  **
        0678: q_reg <= 8'b00111100; // 6   ****
        0679: q_reg <= 8'b11111111; // 7 ********
        0680: q_reg <= 8'b00111100; // 8   ****
        0681: q_reg <= 8'b01100110; // 9  **  **
        0682: q_reg <= 8'b00000000; // a
        0683: q_reg <= 8'b00000000; // b
        0684: q_reg <= 8'b00000000; // c
        0685: q_reg <= 8'b00000000; // d
        0686: q_reg <= 8'b00000000; // e
        0687: q_reg <= 8'b00000000; // f
        // -- code x2b
        0688: q_reg <= 8'b00000000; // 0
        0689: q_reg <= 8'b00000000; // 1
        0690: q_reg <= 8'b00000000; // 2
        0691: q_reg <= 8'b00000000; // 3
        0692: q_reg <= 8'b00000000; // 4
        0693: q_reg <= 8'b00011000; // 5    **
        0694: q_reg <= 8'b00011000; // 6    **
        0695: q_reg <= 8'b01111110; // 7  ******
        0696: q_reg <= 8'b00011000; // 8    **
        0697: q_reg <= 8'b00011000; // 9    **
        0698: q_reg <= 8'b00000000; // a
        0699: q_reg <= 8'b00000000; // b
        0700: q_reg <= 8'b00000000; // c
        0701: q_reg <= 8'b00000000; // d
        0702: q_reg <= 8'b00000000; // e
        0703: q_reg <= 8'b00000000; // f
        // -- code x2c
        0704: q_reg <= 8'b00000000; // 0
        0705: q_reg <= 8'b00000000; // 1
        0706: q_reg <= 8'b00000000; // 2
        0707: q_reg <= 8'b00000000; // 3
        0708: q_reg <= 8'b00000000; // 4
        0709: q_reg <= 8'b00000000; // 5
        0710: q_reg <= 8'b00000000; // 6
        0711: q_reg <= 8'b00000000; // 7
        0712: q_reg <= 8'b00000000; // 8
        0713: q_reg <= 8'b00011000; // 9    **
        0714: q_reg <= 8'b00011000; // a    **
        0715: q_reg <= 8'b00011000; // b    **
        0716: q_reg <= 8'b00110000; // c   **
        0717: q_reg <= 8'b00000000; // d
        0718: q_reg <= 8'b00000000; // e
        0719: q_reg <= 8'b00000000; // f
        // -- code x2d
        0720: q_reg <= 8'b00000000; // 0
        0721: q_reg <= 8'b00000000; // 1
        0722: q_reg <= 8'b00000000; // 2
        0723: q_reg <= 8'b00000000; // 3
        0724: q_reg <= 8'b00000000; // 4
        0725: q_reg <= 8'b00000000; // 5
        0726: q_reg <= 8'b00000000; // 6
        0727: q_reg <= 8'b01111110; // 7  ******
        0728: q_reg <= 8'b00000000; // 8
        0729: q_reg <= 8'b00000000; // 9
        0730: q_reg <= 8'b00000000; // a
        0731: q_reg <= 8'b00000000; // b
        0732: q_reg <= 8'b00000000; // c
        0733: q_reg <= 8'b00000000; // d
        0734: q_reg <= 8'b00000000; // e
        0735: q_reg <= 8'b00000000; // f
        // -- code x2e
        0736: q_reg <= 8'b00000000; // 0
        0737: q_reg <= 8'b00000000; // 1
        0738: q_reg <= 8'b00000000; // 2
        0739: q_reg <= 8'b00000000; // 3
        0740: q_reg <= 8'b00000000; // 4
        0741: q_reg <= 8'b00000000; // 5
        0742: q_reg <= 8'b00000000; // 6
        0743: q_reg <= 8'b00000000; // 7
        0744: q_reg <= 8'b00000000; // 8
        0745: q_reg <= 8'b00000000; // 9
        0746: q_reg <= 8'b00011000; // a    **
        0747: q_reg <= 8'b00011000; // b    **
        0748: q_reg <= 8'b00000000; // c
        0749: q_reg <= 8'b00000000; // d
        0750: q_reg <= 8'b00000000; // e
        0751: q_reg <= 8'b00000000; // f
        // -- code x2f
        0752: q_reg <= 8'b00000000; // 0
        0753: q_reg <= 8'b00000000; // 1
        0754: q_reg <= 8'b00000000; // 2
        0755: q_reg <= 8'b00000000; // 3
        0756: q_reg <= 8'b00000010; // 4       *
        0757: q_reg <= 8'b00000110; // 5      **
        0758: q_reg <= 8'b00001100; // 6     **
        0759: q_reg <= 8'b00011000; // 7    **
        0760: q_reg <= 8'b00110000; // 8   **
        0761: q_reg <= 8'b01100000; // 9  **
        0762: q_reg <= 8'b11000000; // a **
        0763: q_reg <= 8'b10000000; // b *
        0764: q_reg <= 8'b00000000; // c
        0765: q_reg <= 8'b00000000; // d
        0766: q_reg <= 8'b00000000; // e
        0767: q_reg <= 8'b00000000; // f
        // -- 0: code x30
        0768: q_reg <= 8'b00000000; // 0
        0769: q_reg <= 8'b00000000; // 1
        0770: q_reg <= 8'b01111100; // 2  *****
        0771: q_reg <= 8'b11000110; // 3 **   **
        0772: q_reg <= 8'b11000110; // 4 **   **
        0773: q_reg <= 8'b11001110; // 5 **  ***
        0774: q_reg <= 8'b11011110; // 6 ** ****
        0775: q_reg <= 8'b11110110; // 7 **** **
        0776: q_reg <= 8'b11100110; // 8 ***  **
        0777: q_reg <= 8'b11000110; // 9 **   **
        0778: q_reg <= 8'b11000110; // a **   **
        0779: q_reg <= 8'b01111100; // b  *****
        0780: q_reg <= 8'b00000000; // c
        0781: q_reg <= 8'b00000000; // d
        0782: q_reg <= 8'b00000000; // e
        0783: q_reg <= 8'b00000000; // f
        // -- 1: code x31
        0784: q_reg <= 8'b00000000; // 0
        0785: q_reg <= 8'b00000000; // 1
        0786: q_reg <= 8'b00011000; // 2
        0787: q_reg <= 8'b00111000; // 3
        0788: q_reg <= 8'b01111000; // 4    **
        0789: q_reg <= 8'b00011000; // 5   ***
        0790: q_reg <= 8'b00011000; // 6  ****
        0791: q_reg <= 8'b00011000; // 7    **
        0792: q_reg <= 8'b00011000; // 8    **
        0793: q_reg <= 8'b00011000; // 9    **
        0794: q_reg <= 8'b00011000; // a    **
        0795: q_reg <= 8'b01111110; // b    **
        0796: q_reg <= 8'b00000000; // c    **
        0797: q_reg <= 8'b00000000; // d  ******
        0798: q_reg <= 8'b00000000; // e
        0799: q_reg <= 8'b00000000; // f
        // -- 2: code x32
        0800: q_reg <= 8'b00000000; // 0
        0801: q_reg <= 8'b00000000; // 1
        0802: q_reg <= 8'b01111100; // 2  *****
        0803: q_reg <= 8'b11000110; // 3 **   **
        0804: q_reg <= 8'b00000110; // 4      **
        0805: q_reg <= 8'b00001100; // 5     **
        0806: q_reg <= 8'b00011000; // 6    **
        0807: q_reg <= 8'b00110000; // 7   **
        0808: q_reg <= 8'b01100000; // 8  **
        0809: q_reg <= 8'b11000000; // 9 **
        0810: q_reg <= 8'b11000110; // a **   **
        0811: q_reg <= 8'b11111110; // b *******
        0812: q_reg <= 8'b00000000; // c
        0813: q_reg <= 8'b00000000; // d
        0814: q_reg <= 8'b00000000; // e
        0815: q_reg <= 8'b00000000; // f
        // -- 3: code x33
        0816: q_reg <= 8'b00000000; // 0
        0817: q_reg <= 8'b00000000; // 1
        0818: q_reg <= 8'b01111100; // 2  *****
        0819: q_reg <= 8'b11000110; // 3 **   **
        0820: q_reg <= 8'b00000110; // 4      **
        0821: q_reg <= 8'b00000110; // 5      **
        0822: q_reg <= 8'b00111100; // 6   ****
        0823: q_reg <= 8'b00000110; // 7      **
        0824: q_reg <= 8'b00000110; // 8      **
        0825: q_reg <= 8'b00000110; // 9      **
        0826: q_reg <= 8'b11000110; // a **   **
        0827: q_reg <= 8'b01111100; // b  *****
        0828: q_reg <= 8'b00000000; // c
        0829: q_reg <= 8'b00000000; // d
        0830: q_reg <= 8'b00000000; // e
        0831: q_reg <= 8'b00000000; // f
        // -- 4: code x34
        0832: q_reg <= 8'b00000000; // 0
        0833: q_reg <= 8'b00000000; // 1
        0834: q_reg <= 8'b00001100; // 2     **
        0835: q_reg <= 8'b00011100; // 3    ***
        0836: q_reg <= 8'b00111100; // 4   ****
        0837: q_reg <= 8'b01101100; // 5  ** **
        0838: q_reg <= 8'b11001100; // 6 **  **
        0839: q_reg <= 8'b11111110; // 7 *******
        0840: q_reg <= 8'b00001100; // 8     **
        0841: q_reg <= 8'b00001100; // 9     **
        0842: q_reg <= 8'b00001100; // a     **
        0843: q_reg <= 8'b00011110; // b    ****
        0844: q_reg <= 8'b00000000; // c
        0845: q_reg <= 8'b00000000; // d
        0846: q_reg <= 8'b00000000; // e
        0847: q_reg <= 8'b00000000; // f
        // -- code x35
        0848: q_reg <= 8'b00000000; // 0
        0849: q_reg <= 8'b00000000; // 1
        0850: q_reg <= 8'b11111110; // 2 *******
        0851: q_reg <= 8'b11000000; // 3 **
        0852: q_reg <= 8'b11000000; // 4 **
        0853: q_reg <= 8'b11000000; // 5 **
        0854: q_reg <= 8'b11111100; // 6 ******
        0855: q_reg <= 8'b00000110; // 7      **
        0856: q_reg <= 8'b00000110; // 8      **
        0857: q_reg <= 8'b00000110; // 9      **
        0858: q_reg <= 8'b11000110; // a **   **
        0859: q_reg <= 8'b01111100; // b  *****
        0860: q_reg <= 8'b00000000; // c
        0861: q_reg <= 8'b00000000; // d
        0862: q_reg <= 8'b00000000; // e
        0863: q_reg <= 8'b00000000; // f
        // -- code x36
        0864: q_reg <= 8'b00000000; // 0
        0865: q_reg <= 8'b00000000; // 1
        0866: q_reg <= 8'b00111000; // 2   ***
        0867: q_reg <= 8'b01100000; // 3  **
        0868: q_reg <= 8'b11000000; // 4 **
        0869: q_reg <= 8'b11000000; // 5 **
        0870: q_reg <= 8'b11111100; // 6 ******
        0871: q_reg <= 8'b11000110; // 7 **   **
        0872: q_reg <= 8'b11000110; // 8 **   **
        0873: q_reg <= 8'b11000110; // 9 **   **
        0874: q_reg <= 8'b11000110; // a **   **
        0875: q_reg <= 8'b01111100; // b  *****
        0876: q_reg <= 8'b00000000; // c
        0877: q_reg <= 8'b00000000; // d
        0878: q_reg <= 8'b00000000; // e
        0879: q_reg <= 8'b00000000; // f
        // -- code x37
        0880: q_reg <= 8'b00000000; // 0
        0881: q_reg <= 8'b00000000; // 1
        0882: q_reg <= 8'b11111110; // 2 *******
        0883: q_reg <= 8'b11000110; // 3 **   **
        0884: q_reg <= 8'b00000110; // 4      **
        0885: q_reg <= 8'b00000110; // 5      **
        0886: q_reg <= 8'b00001100; // 6     **
        0887: q_reg <= 8'b00011000; // 7    **
        0888: q_reg <= 8'b00110000; // 8   **
        0889: q_reg <= 8'b00110000; // 9   **
        0890: q_reg <= 8'b00110000; // a   **
        0891: q_reg <= 8'b00110000; // b   **
        0892: q_reg <= 8'b00000000; // c
        0893: q_reg <= 8'b00000000; // d
        0894: q_reg <= 8'b00000000; // e
        0895: q_reg <= 8'b00000000; // f
        // -- code x38
        0896: q_reg <= 8'b00000000; // 0
        0897: q_reg <= 8'b00000000; // 1
        0898: q_reg <= 8'b01111100; // 2  *****
        0899: q_reg <= 8'b11000110; // 3 **   **
        0900: q_reg <= 8'b11000110; // 4 **   **
        0901: q_reg <= 8'b11000110; // 5 **   **
        0902: q_reg <= 8'b01111100; // 6  *****
        0903: q_reg <= 8'b11000110; // 7 **   **
        0904: q_reg <= 8'b11000110; // 8 **   **
        0905: q_reg <= 8'b11000110; // 9 **   **
        0906: q_reg <= 8'b11000110; // a **   **
        0907: q_reg <= 8'b01111100; // b  *****
        0908: q_reg <= 8'b00000000; // c
        0909: q_reg <= 8'b00000000; // d
        0910: q_reg <= 8'b00000000; // e
        0911: q_reg <= 8'b00000000; // f
        // -- code x39
        0912: q_reg <= 8'b00000000; // 0
        0913: q_reg <= 8'b00000000; // 1
        0914: q_reg <= 8'b01111100; // 2  *****
        0915: q_reg <= 8'b11000110; // 3 **   **
        0916: q_reg <= 8'b11000110; // 4 **   **
        0917: q_reg <= 8'b11000110; // 5 **   **
        0918: q_reg <= 8'b01111110; // 6  ******
        0919: q_reg <= 8'b00000110; // 7      **
        0920: q_reg <= 8'b00000110; // 8      **
        0921: q_reg <= 8'b00000110; // 9      **
        0922: q_reg <= 8'b00001100; // a     **
        0923: q_reg <= 8'b01111000; // b  ****
        0924: q_reg <= 8'b00000000; // c
        0925: q_reg <= 8'b00000000; // d
        0926: q_reg <= 8'b00000000; // e
        0927: q_reg <= 8'b00000000; // f
        // -- code x3a
        0928: q_reg <= 8'b00000000; // 0
        0929: q_reg <= 8'b00000000; // 1
        0930: q_reg <= 8'b00000000; // 2
        0931: q_reg <= 8'b00000000; // 3
        0932: q_reg <= 8'b00011000; // 4    **
        0933: q_reg <= 8'b00011000; // 5    **
        0934: q_reg <= 8'b00000000; // 6
        0935: q_reg <= 8'b00000000; // 7
        0936: q_reg <= 8'b00000000; // 8
        0937: q_reg <= 8'b00011000; // 9    **
        0938: q_reg <= 8'b00011000; // a    **
        0939: q_reg <= 8'b00000000; // b
        0940: q_reg <= 8'b00000000; // c
        0941: q_reg <= 8'b00000000; // d
        0942: q_reg <= 8'b00000000; // e
        0943: q_reg <= 8'b00000000; // f
        // -- code x3b
        0944: q_reg <= 8'b00000000; // 0
        0945: q_reg <= 8'b00000000; // 1
        0946: q_reg <= 8'b00000000; // 2
        0947: q_reg <= 8'b00000000; // 3
        0948: q_reg <= 8'b00011000; // 4    **
        0949: q_reg <= 8'b00011000; // 5    **
        0950: q_reg <= 8'b00000000; // 6
        0951: q_reg <= 8'b00000000; // 7
        0952: q_reg <= 8'b00000000; // 8
        0953: q_reg <= 8'b00011000; // 9    **
        0954: q_reg <= 8'b00011000; // a    **
        0955: q_reg <= 8'b00110000; // b   **
        0956: q_reg <= 8'b00000000; // c
        0957: q_reg <= 8'b00000000; // d
        0958: q_reg <= 8'b00000000; // e
        0959: q_reg <= 8'b00000000; // f
        // -- code x3c
        0960: q_reg <= 8'b00000000; // 0
        0961: q_reg <= 8'b00000000; // 1
        0962: q_reg <= 8'b00000000; // 2
        0963: q_reg <= 8'b00000110; // 3      **
        0964: q_reg <= 8'b00001100; // 4     **
        0965: q_reg <= 8'b00011000; // 5    **
        0966: q_reg <= 8'b00110000; // 6   **
        0967: q_reg <= 8'b01100000; // 7  **
        0968: q_reg <= 8'b00110000; // 8   **
        0969: q_reg <= 8'b00011000; // 9    **
        0970: q_reg <= 8'b00001100; // a     **
        0971: q_reg <= 8'b00000110; // b      **
        0972: q_reg <= 8'b00000000; // c
        0973: q_reg <= 8'b00000000; // d
        0974: q_reg <= 8'b00000000; // e
        0975: q_reg <= 8'b00000000; // f
        // -- code x3d
        0976: q_reg <= 8'b00000000; // 0
        0977: q_reg <= 8'b00000000; // 1
        0978: q_reg <= 8'b00000000; // 2
        0979: q_reg <= 8'b00000000; // 3
        0980: q_reg <= 8'b00000000; // 4
        0981: q_reg <= 8'b01111110; // 5  ******
        0982: q_reg <= 8'b00000000; // 6
        0983: q_reg <= 8'b00000000; // 7
        0984: q_reg <= 8'b01111110; // 8  ******
        0985: q_reg <= 8'b00000000; // 9
        0986: q_reg <= 8'b00000000; // a
        0987: q_reg <= 8'b00000000; // b
        0988: q_reg <= 8'b00000000; // c
        0989: q_reg <= 8'b00000000; // d
        0990: q_reg <= 8'b00000000; // e
        0991: q_reg <= 8'b00000000; // f
        // -- code x3e
        0992: q_reg <= 8'b00000000; // 0
        0993: q_reg <= 8'b00000000; // 1
        0994: q_reg <= 8'b00000000; // 2
        0995: q_reg <= 8'b01100000; // 3  **
        0996: q_reg <= 8'b00110000; // 4   **
        0997: q_reg <= 8'b00011000; // 5    **
        0998: q_reg <= 8'b00001100; // 6     **
        0999: q_reg <= 8'b00000110; // 7      **
        1000: q_reg <= 8'b00001100; // 8     **
        1001: q_reg <= 8'b00011000; // 9    **
        1002: q_reg <= 8'b00110000; // a   **
        1003: q_reg <= 8'b01100000; // b  **
        1004: q_reg <= 8'b00000000; // c
        1005: q_reg <= 8'b00000000; // d
        1006: q_reg <= 8'b00000000; // e
        1007: q_reg <= 8'b00000000; // f
        // -- code x3f
        1008: q_reg <= 8'b00000000; // 0
        1009: q_reg <= 8'b00000000; // 1
        1010: q_reg <= 8'b01111100; // 2  *****
        1011: q_reg <= 8'b11000110; // 3 **   **
        1012: q_reg <= 8'b11000110; // 4 **   **
        1013: q_reg <= 8'b00001100; // 5     **
        1014: q_reg <= 8'b00011000; // 6    **
        1015: q_reg <= 8'b00011000; // 7    **
        1016: q_reg <= 8'b00011000; // 8    **
        1017: q_reg <= 8'b00000000; // 9
        1018: q_reg <= 8'b00011000; // a    **
        1019: q_reg <= 8'b00011000; // b    **
        1020: q_reg <= 8'b00000000; // c
        1021: q_reg <= 8'b00000000; // d
        1022: q_reg <= 8'b00000000; // e
        1023: q_reg <= 8'b00000000; // f
        // -- code x40
        1024: q_reg <= 8'b00000000; // 0
        1025: q_reg <= 8'b00000000; // 1
        1026: q_reg <= 8'b01111100; // 2  *****
        1027: q_reg <= 8'b11000110; // 3 **   **
        1028: q_reg <= 8'b11000110; // 4 **   **
        1029: q_reg <= 8'b11000110; // 5 **   **
        1030: q_reg <= 8'b11011110; // 6 ** ****
        1031: q_reg <= 8'b11011110; // 7 ** ****
        1032: q_reg <= 8'b11011110; // 8 ** ****
        1033: q_reg <= 8'b11011100; // 9 ** ***
        1034: q_reg <= 8'b11000000; // a **
        1035: q_reg <= 8'b01111100; // b  *****
        1036: q_reg <= 8'b00000000; // c
        1037: q_reg <= 8'b00000000; // d
        1038: q_reg <= 8'b00000000; // e
        1039: q_reg <= 8'b00000000; // f
        // -- A: code x41
        1040: q_reg <= 8'b00000000; // 0
        1041: q_reg <= 8'b00000000; // 1
        1042: q_reg <= 8'b00010000; // 2    *
        1043: q_reg <= 8'b00111000; // 3   ***
        1044: q_reg <= 8'b01101100; // 4  ** **
        1045: q_reg <= 8'b11000110; // 5 **   **
        1046: q_reg <= 8'b11000110; // 6 **   **
        1047: q_reg <= 8'b11111110; // 7 *******
        1048: q_reg <= 8'b11000110; // 8 **   **
        1049: q_reg <= 8'b11000110; // 9 **   **
        1050: q_reg <= 8'b11000110; // a **   **
        1051: q_reg <= 8'b11000110; // b **   **
        1052: q_reg <= 8'b00000000; // c
        1053: q_reg <= 8'b00000000; // d
        1054: q_reg <= 8'b00000000; // e
        1055: q_reg <= 8'b00000000; // f
        // -- B: code x42
        1056: q_reg <= 8'b00000000; // 0
        1057: q_reg <= 8'b00000000; // 1
        1058: q_reg <= 8'b11111100; // 2 ******
        1059: q_reg <= 8'b01100110; // 3  **  **
        1060: q_reg <= 8'b01100110; // 4  **  **
        1061: q_reg <= 8'b01100110; // 5  **  **
        1062: q_reg <= 8'b01111100; // 6  *****
        1063: q_reg <= 8'b01100110; // 7  **  **
        1064: q_reg <= 8'b01100110; // 8  **  **
        1065: q_reg <= 8'b01100110; // 9  **  **
        1066: q_reg <= 8'b01100110; // a  **  **
        1067: q_reg <= 8'b11111100; // b ******
        1068: q_reg <= 8'b00000000; // c
        1069: q_reg <= 8'b00000000; // d
        1070: q_reg <= 8'b00000000; // e
        1071: q_reg <= 8'b00000000; // f
        // -- C: code x43
        1072: q_reg <= 8'b00000000; // 0
        1073: q_reg <= 8'b00000000; // 1
        1074: q_reg <= 8'b00111100; // 2   ****
        1075: q_reg <= 8'b01100110; // 3  **  **
        1076: q_reg <= 8'b11000010; // 4 **    *
        1077: q_reg <= 8'b11000000; // 5 **
        1078: q_reg <= 8'b11000000; // 6 **
        1079: q_reg <= 8'b11000000; // 7 **
        1080: q_reg <= 8'b11000000; // 8 **
        1081: q_reg <= 8'b11000010; // 9 **    *
        1082: q_reg <= 8'b01100110; // a  **  **
        1083: q_reg <= 8'b00111100; // b   ****
        1084: q_reg <= 8'b00000000; // c
        1085: q_reg <= 8'b00000000; // d
        1086: q_reg <= 8'b00000000; // e
        1087: q_reg <= 8'b00000000; // f
        // -- D: code x44
        1088: q_reg <= 8'b00000000; // 0
        1089: q_reg <= 8'b00000000; // 1
        1090: q_reg <= 8'b11111000; // 2 *****
        1091: q_reg <= 8'b01101100; // 3  ** **
        1092: q_reg <= 8'b01100110; // 4  **  **
        1093: q_reg <= 8'b01100110; // 5  **  **
        1094: q_reg <= 8'b01100110; // 6  **  **
        1095: q_reg <= 8'b01100110; // 7  **  **
        1096: q_reg <= 8'b01100110; // 8  **  **
        1097: q_reg <= 8'b01100110; // 9  **  **
        1098: q_reg <= 8'b01101100; // a  ** **
        1099: q_reg <= 8'b11111000; // b *****
        1100: q_reg <= 8'b00000000; // c
        1101: q_reg <= 8'b00000000; // d
        1102: q_reg <= 8'b00000000; // e
        1103: q_reg <= 8'b00000000; // f
        // -- code x45
        1104: q_reg <= 8'b00000000; // 0
        1105: q_reg <= 8'b00000000; // 1
        1106: q_reg <= 8'b11111110; // 2 *******
        1107: q_reg <= 8'b01100110; // 3  **  **
        1108: q_reg <= 8'b01100010; // 4  **   *
        1109: q_reg <= 8'b01101000; // 5  ** *
        1110: q_reg <= 8'b01111000; // 6  ****
        1111: q_reg <= 8'b01101000; // 7  ** *
        1112: q_reg <= 8'b01100000; // 8  **
        1113: q_reg <= 8'b01100010; // 9  **   *
        1114: q_reg <= 8'b01100110; // a  **  **
        1115: q_reg <= 8'b11111110; // b *******
        1116: q_reg <= 8'b00000000; // c
        1117: q_reg <= 8'b00000000; // d
        1118: q_reg <= 8'b00000000; // e
        1119: q_reg <= 8'b00000000; // f
        // -- code x46
        1120: q_reg <= 8'b00000000; // 0
        1121: q_reg <= 8'b00000000; // 1
        1122: q_reg <= 8'b11111110; // 2 *******
        1123: q_reg <= 8'b01100110; // 3  **  **
        1124: q_reg <= 8'b01100010; // 4  **   *
        1125: q_reg <= 8'b01101000; // 5  ** *
        1126: q_reg <= 8'b01111000; // 6  ****
        1127: q_reg <= 8'b01101000; // 7  ** *
        1128: q_reg <= 8'b01100000; // 8  **
        1129: q_reg <= 8'b01100000; // 9  **
        1130: q_reg <= 8'b01100000; // a  **
        1131: q_reg <= 8'b11110000; // b ****
        1132: q_reg <= 8'b00000000; // c
        1133: q_reg <= 8'b00000000; // d
        1134: q_reg <= 8'b00000000; // e
        1135: q_reg <= 8'b00000000; // f
        // -- code x47
        1136: q_reg <= 8'b00000000; // 0
        1137: q_reg <= 8'b00000000; // 1
        1138: q_reg <= 8'b00111100; // 2   ****
        1139: q_reg <= 8'b01100110; // 3  **  **
        1140: q_reg <= 8'b11000010; // 4 **    *
        1141: q_reg <= 8'b11000000; // 5 **
        1142: q_reg <= 8'b11000000; // 6 **
        1143: q_reg <= 8'b11011110; // 7 ** ****
        1144: q_reg <= 8'b11000110; // 8 **   **
        1145: q_reg <= 8'b11000110; // 9 **   **
        1146: q_reg <= 8'b01100110; // a  **  **
        1147: q_reg <= 8'b00111010; // b   *** *
        1148: q_reg <= 8'b00000000; // c
        1149: q_reg <= 8'b00000000; // d
        1150: q_reg <= 8'b00000000; // e
        1151: q_reg <= 8'b00000000; // f
        // -- H: code x48
        1152: q_reg <= 8'b00000000; // 0
        1153: q_reg <= 8'b00000000; // 1
        1154: q_reg <= 8'b11000110; // 2 **   **
        1155: q_reg <= 8'b11000110; // 3 **   **
        1156: q_reg <= 8'b11000110; // 4 **   **
        1157: q_reg <= 8'b11000110; // 5 **   **
        1158: q_reg <= 8'b11111110; // 6 *******
        1159: q_reg <= 8'b11000110; // 7 **   **
        1160: q_reg <= 8'b11000110; // 8 **   **
        1161: q_reg <= 8'b11000110; // 9 **   **
        1162: q_reg <= 8'b11000110; // a **   **
        1163: q_reg <= 8'b11000110; // b **   **
        1164: q_reg <= 8'b00000000; // c
        1165: q_reg <= 8'b00000000; // d
        1166: q_reg <= 8'b00000000; // e
        1167: q_reg <= 8'b00000000; // f
        // -- I: code x49
        1168: q_reg <= 8'b00000000; // 0
        1169: q_reg <= 8'b00000000; // 1
        1170: q_reg <= 8'b00111100; // 2   ****
        1171: q_reg <= 8'b00011000; // 3    **
        1172: q_reg <= 8'b00011000; // 4    **
        1173: q_reg <= 8'b00011000; // 5    **
        1174: q_reg <= 8'b00011000; // 6    **
        1175: q_reg <= 8'b00011000; // 7    **
        1176: q_reg <= 8'b00011000; // 8    **
        1177: q_reg <= 8'b00011000; // 9    **
        1178: q_reg <= 8'b00011000; // a    **
        1179: q_reg <= 8'b00111100; // b   ****
        1180: q_reg <= 8'b00000000; // c
        1181: q_reg <= 8'b00000000; // d
        1182: q_reg <= 8'b00000000; // e
        1183: q_reg <= 8'b00000000; // f
        // -- J: code x4a
        1184: q_reg <= 8'b00000000; // 0
        1185: q_reg <= 8'b00000000; // 1
        1186: q_reg <= 8'b00011110; // 2    ****
        1187: q_reg <= 8'b00001100; // 3     **
        1188: q_reg <= 8'b00001100; // 4     **
        1189: q_reg <= 8'b00001100; // 5     **
        1190: q_reg <= 8'b00001100; // 6     **
        1191: q_reg <= 8'b00001100; // 7     **
        1192: q_reg <= 8'b11001100; // 8 **  **
        1193: q_reg <= 8'b11001100; // 9 **  **
        1194: q_reg <= 8'b11001100; // a **  **
        1195: q_reg <= 8'b01111000; // b  ****
        1196: q_reg <= 8'b00000000; // c
        1197: q_reg <= 8'b00000000; // d
        1198: q_reg <= 8'b00000000; // e
        1199: q_reg <= 8'b00000000; // f
        // -- K: code x4b
        1200: q_reg <= 8'b00000000; // 0
        1201: q_reg <= 8'b00000000; // 1
        1202: q_reg <= 8'b11100110; // 2 ***  **
        1203: q_reg <= 8'b01100110; // 3  **  **
        1204: q_reg <= 8'b01100110; // 4  **  **
        1205: q_reg <= 8'b01101100; // 5  ** **
        1206: q_reg <= 8'b01111000; // 6  ****
        1207: q_reg <= 8'b01111000; // 7  ****
        1208: q_reg <= 8'b01101100; // 8  ** **
        1209: q_reg <= 8'b01100110; // 9  **  **
        1210: q_reg <= 8'b01100110; // a  **  **
        1211: q_reg <= 8'b11100110; // b ***  **
        1212: q_reg <= 8'b00000000; // c
        1213: q_reg <= 8'b00000000; // d
        1214: q_reg <= 8'b00000000; // e
        1215: q_reg <= 8'b00000000; // f
        // -- L: code x4c
        1216: q_reg <= 8'b00000000; // 0
        1217: q_reg <= 8'b00000000; // 1
        1218: q_reg <= 8'b11110000; // 2 ****
        1219: q_reg <= 8'b01100000; // 3  **
        1220: q_reg <= 8'b01100000; // 4  **
        1221: q_reg <= 8'b01100000; // 5  **
        1222: q_reg <= 8'b01100000; // 6  **
        1223: q_reg <= 8'b01100000; // 7  **
        1224: q_reg <= 8'b01100000; // 8  **
        1225: q_reg <= 8'b01100010; // 9  **   *
        1226: q_reg <= 8'b01100110; // a  **  **
        1227: q_reg <= 8'b11111110; // b *******
        1228: q_reg <= 8'b00000000; // c
        1229: q_reg <= 8'b00000000; // d
        1230: q_reg <= 8'b00000000; // e
        1231: q_reg <= 8'b00000000; // f
        // -- M: code x4d
        1232: q_reg <= 8'b00000000; // 0
        1233: q_reg <= 8'b00000000; // 1
        1234: q_reg <= 8'b11000011; // 2 **    **
        1235: q_reg <= 8'b11100111; // 3 ***  ***
        1236: q_reg <= 8'b11111111; // 4 ********
        1237: q_reg <= 8'b11111111; // 5 ********
        1238: q_reg <= 8'b11011011; // 6 ** ** **
        1239: q_reg <= 8'b11000011; // 7 **    **
        1240: q_reg <= 8'b11000011; // 8 **    **
        1241: q_reg <= 8'b11000011; // 9 **    **
        1242: q_reg <= 8'b11000011; // a **    **
        1243: q_reg <= 8'b11000011; // b **    **
        1244: q_reg <= 8'b00000000; // c
        1245: q_reg <= 8'b00000000; // d
        1246: q_reg <= 8'b00000000; // e
        1247: q_reg <= 8'b00000000; // f
        // -- N: code x4e
        1248: q_reg <= 8'b00000000; // 0
        1249: q_reg <= 8'b00000000; // 1
        1250: q_reg <= 8'b11000110; // 2 **   **
        1251: q_reg <= 8'b11100110; // 3 ***  **
        1252: q_reg <= 8'b11110110; // 4 **** **
        1253: q_reg <= 8'b11111110; // 5 *******
        1254: q_reg <= 8'b11011110; // 6 ** ****
        1255: q_reg <= 8'b11001110; // 7 **  ***
        1256: q_reg <= 8'b11000110; // 8 **   **
        1257: q_reg <= 8'b11000110; // 9 **   **
        1258: q_reg <= 8'b11000110; // a **   **
        1259: q_reg <= 8'b11000110; // b **   **
        1260: q_reg <= 8'b00000000; // c
        1261: q_reg <= 8'b00000000; // d
        1262: q_reg <= 8'b00000000; // e
        1263: q_reg <= 8'b00000000; // f
        // -- O: code x4f
        1264: q_reg <= 8'b00000000; // 0
        1265: q_reg <= 8'b00000000; // 1
        1266: q_reg <= 8'b01111100; // 2  *****
        1267: q_reg <= 8'b11000110; // 3 **   **
        1268: q_reg <= 8'b11000110; // 4 **   **
        1269: q_reg <= 8'b11000110; // 5 **   **
        1270: q_reg <= 8'b11000110; // 6 **   **
        1271: q_reg <= 8'b11000110; // 7 **   **
        1272: q_reg <= 8'b11000110; // 8 **   **
        1273: q_reg <= 8'b11000110; // 9 **   **
        1274: q_reg <= 8'b11000110; // a **   **
        1275: q_reg <= 8'b01111100; // b  *****
        1276: q_reg <= 8'b00000000; // c
        1277: q_reg <= 8'b00000000; // d
        1278: q_reg <= 8'b00000000; // e
        1279: q_reg <= 8'b00000000; // f
        // -- P: code x50
        1280: q_reg <= 8'b00000000; // 0
        1281: q_reg <= 8'b00000000; // 1
        1282: q_reg <= 8'b11111100; // 2 ******
        1283: q_reg <= 8'b01100110; // 3  **  **
        1284: q_reg <= 8'b01100110; // 4  **  **
        1285: q_reg <= 8'b01100110; // 5  **  **
        1286: q_reg <= 8'b01111100; // 6  *****
        1287: q_reg <= 8'b01100000; // 7  **
        1288: q_reg <= 8'b01100000; // 8  **
        1289: q_reg <= 8'b01100000; // 9  **
        1290: q_reg <= 8'b01100000; // a  **
        1291: q_reg <= 8'b11110000; // b ****
        1292: q_reg <= 8'b00000000; // c
        1293: q_reg <= 8'b00000000; // d
        1294: q_reg <= 8'b00000000; // e
        1295: q_reg <= 8'b00000000; // f
        // -- Q: code x510
        1296: q_reg <= 8'b00000000; // 0
        1297: q_reg <= 8'b00000000; // 1
        1298: q_reg <= 8'b01111100; // 2  *****
        1299: q_reg <= 8'b11000110; // 3 **   **
        1300: q_reg <= 8'b11000110; // 4 **   **
        1301: q_reg <= 8'b11000110; // 5 **   **
        1302: q_reg <= 8'b11000110; // 6 **   **
        1303: q_reg <= 8'b11000110; // 7 **   **
        1304: q_reg <= 8'b11000110; // 8 **   **
        1305: q_reg <= 8'b11010110; // 9 ** * **
        1306: q_reg <= 8'b11011110; // a ** ****
        1307: q_reg <= 8'b01111100; // b  *****
        1308: q_reg <= 8'b00001100; // c     **
        1309: q_reg <= 8'b00001110; // d     ***
        1310: q_reg <= 8'b00000000; // e
        1311: q_reg <= 8'b00000000; // f
        // -- code x52
        1312: q_reg <= 8'b00000000; // 0
        1313: q_reg <= 8'b00000000; // 1
        1314: q_reg <= 8'b11111100; // 2 ******
        1315: q_reg <= 8'b01100110; // 3  **  **
        1316: q_reg <= 8'b01100110; // 4  **  **
        1317: q_reg <= 8'b01100110; // 5  **  **
        1318: q_reg <= 8'b01111100; // 6  *****
        1319: q_reg <= 8'b01101100; // 7  ** **
        1320: q_reg <= 8'b01100110; // 8  **  **
        1321: q_reg <= 8'b01100110; // 9  **  **
        1322: q_reg <= 8'b01100110; // a  **  **
        1323: q_reg <= 8'b11100110; // b ***  **
        1324: q_reg <= 8'b00000000; // c
        1325: q_reg <= 8'b00000000; // d
        1326: q_reg <= 8'b00000000; // e
        1327: q_reg <= 8'b00000000; // f
        // -- code x53
        1328: q_reg <= 8'b00000000; // 0
        1329: q_reg <= 8'b00000000; // 1
        1330: q_reg <= 8'b01111100; // 2  *****
        1331: q_reg <= 8'b11000110; // 3 **   **
        1332: q_reg <= 8'b11000110; // 4 **   **
        1333: q_reg <= 8'b01100000; // 5  **
        1334: q_reg <= 8'b00111000; // 6   ***
        1335: q_reg <= 8'b00001100; // 7     **
        1336: q_reg <= 8'b00000110; // 8      **
        1337: q_reg <= 8'b11000110; // 9 **   **
        1338: q_reg <= 8'b11000110; // a **   **
        1339: q_reg <= 8'b01111100; // b  *****
        1340: q_reg <= 8'b00000000; // c
        1341: q_reg <= 8'b00000000; // d
        1342: q_reg <= 8'b00000000; // e
        1343: q_reg <= 8'b00000000; // f
        // -- code x54
        1344: q_reg <= 8'b00000000; // 0
        1345: q_reg <= 8'b00000000; // 1
        1346: q_reg <= 8'b11111111; // 2 ********
        1347: q_reg <= 8'b11011011; // 3 ** ** **
        1348: q_reg <= 8'b10011001; // 4 *  **  *
        1349: q_reg <= 8'b00011000; // 5    **
        1350: q_reg <= 8'b00011000; // 6    **
        1351: q_reg <= 8'b00011000; // 7    **
        1352: q_reg <= 8'b00011000; // 8    **
        1353: q_reg <= 8'b00011000; // 9    **
        1354: q_reg <= 8'b00011000; // a    **
        1355: q_reg <= 8'b00111100; // b   ****
        1356: q_reg <= 8'b00000000; // c
        1357: q_reg <= 8'b00000000; // d
        1358: q_reg <= 8'b00000000; // e
        1359: q_reg <= 8'b00000000; // f
        // -- code x55
        1360: q_reg <= 8'b00000000; // 0
        1361: q_reg <= 8'b00000000; // 1
        1362: q_reg <= 8'b11000110; // 2 **   **
        1363: q_reg <= 8'b11000110; // 3 **   **
        1364: q_reg <= 8'b11000110; // 4 **   **
        1365: q_reg <= 8'b11000110; // 5 **   **
        1366: q_reg <= 8'b11000110; // 6 **   **
        1367: q_reg <= 8'b11000110; // 7 **   **
        1368: q_reg <= 8'b11000110; // 8 **   **
        1369: q_reg <= 8'b11000110; // 9 **   **
        1370: q_reg <= 8'b11000110; // a **   **
        1371: q_reg <= 8'b01111100; // b  *****
        1372: q_reg <= 8'b00000000; // c
        1373: q_reg <= 8'b00000000; // d
        1374: q_reg <= 8'b00000000; // e
        1375: q_reg <= 8'b00000000; // f
        // -- code x56
        1376: q_reg <= 8'b00000000; // 0
        1377: q_reg <= 8'b00000000; // 1
        1378: q_reg <= 8'b11000011; // 2 **    **
        1379: q_reg <= 8'b11000011; // 3 **    **
        1380: q_reg <= 8'b11000011; // 4 **    **
        1381: q_reg <= 8'b11000011; // 5 **    **
        1382: q_reg <= 8'b11000011; // 6 **    **
        1383: q_reg <= 8'b11000011; // 7 **    **
        1384: q_reg <= 8'b11000011; // 8 **    **
        1385: q_reg <= 8'b01100110; // 9  **  **
        1386: q_reg <= 8'b00111100; // a   ****
        1387: q_reg <= 8'b00011000; // b    **
        1388: q_reg <= 8'b00000000; // c
        1389: q_reg <= 8'b00000000; // d
        1390: q_reg <= 8'b00000000; // e
        1391: q_reg <= 8'b00000000; // f
        // -- code x57
        1392: q_reg <= 8'b00000000; // 0
        1393: q_reg <= 8'b00000000; // 1
        1394: q_reg <= 8'b11000011; // 2 **    **
        1395: q_reg <= 8'b11000011; // 3 **    **
        1396: q_reg <= 8'b11000011; // 4 **    **
        1397: q_reg <= 8'b11000011; // 5 **    **
        1398: q_reg <= 8'b11000011; // 6 **    **
        1399: q_reg <= 8'b11011011; // 7 ** ** **
        1400: q_reg <= 8'b11011011; // 8 ** ** **
        1401: q_reg <= 8'b11111111; // 9 ********
        1402: q_reg <= 8'b01100110; // a  **  **
        1403: q_reg <= 8'b01100110; // b  **  **
        1404: q_reg <= 8'b00000000; // c
        1405: q_reg <= 8'b00000000; // d
        1406: q_reg <= 8'b00000000; // e
        1407: q_reg <= 8'b00000000; // f
        // -- code x58
        1408: q_reg <= 8'b00000000; // 0
        1409: q_reg <= 8'b00000000; // 1
        1410: q_reg <= 8'b11000011; // 2 **    **
        1411: q_reg <= 8'b11000011; // 3 **    **
        1412: q_reg <= 8'b01100110; // 4  **  **
        1413: q_reg <= 8'b00111100; // 5   ****
        1414: q_reg <= 8'b00011000; // 6    **
        1415: q_reg <= 8'b00011000; // 7    **
        1416: q_reg <= 8'b00111100; // 8   ****
        1417: q_reg <= 8'b01100110; // 9  **  **
        1418: q_reg <= 8'b11000011; // a **    **
        1419: q_reg <= 8'b11000011; // b **    **
        1420: q_reg <= 8'b00000000; // c
        1421: q_reg <= 8'b00000000; // d
        1422: q_reg <= 8'b00000000; // e
        1423: q_reg <= 8'b00000000; // f
        // -- code x59
        1424: q_reg <= 8'b00000000; // 0
        1425: q_reg <= 8'b00000000; // 1
        1426: q_reg <= 8'b11000011; // 2 **    **
        1427: q_reg <= 8'b11000011; // 3 **    **
        1428: q_reg <= 8'b11000011; // 4 **    **
        1429: q_reg <= 8'b01100110; // 5  **  **
        1430: q_reg <= 8'b00111100; // 6   ****
        1431: q_reg <= 8'b00011000; // 7    **
        1432: q_reg <= 8'b00011000; // 8    **
        1433: q_reg <= 8'b00011000; // 9    **
        1434: q_reg <= 8'b00011000; // a    **
        1435: q_reg <= 8'b00111100; // b   ****
        1436: q_reg <= 8'b00000000; // c
        1437: q_reg <= 8'b00000000; // d
        1438: q_reg <= 8'b00000000; // e
        1439: q_reg <= 8'b00000000; // f
        // -- code x5a
        1440: q_reg <= 8'b00000000; // 0
        1441: q_reg <= 8'b00000000; // 1
        1442: q_reg <= 8'b11111111; // 2 ********
        1443: q_reg <= 8'b11000011; // 3 **    **
        1444: q_reg <= 8'b10000110; // 4 *    **
        1445: q_reg <= 8'b00001100; // 5     **
        1446: q_reg <= 8'b00011000; // 6    **
        1447: q_reg <= 8'b00110000; // 7   **
        1448: q_reg <= 8'b01100000; // 8  **
        1449: q_reg <= 8'b11000001; // 9 **     *
        1450: q_reg <= 8'b11000011; // a **    **
        1451: q_reg <= 8'b11111111; // b ********
        1452: q_reg <= 8'b00000000; // c
        1453: q_reg <= 8'b00000000; // d
        1454: q_reg <= 8'b00000000; // e
        1455: q_reg <= 8'b00000000; // f
        // -- code x5b
        1456: q_reg <= 8'b00000000; // 0
        1457: q_reg <= 8'b00000000; // 1
        1458: q_reg <= 8'b00111100; // 2   ****
        1459: q_reg <= 8'b00110000; // 3   **
        1460: q_reg <= 8'b00110000; // 4   **
        1461: q_reg <= 8'b00110000; // 5   **
        1462: q_reg <= 8'b00110000; // 6   **
        1463: q_reg <= 8'b00110000; // 7   **
        1464: q_reg <= 8'b00110000; // 8   **
        1465: q_reg <= 8'b00110000; // 9   **
        1466: q_reg <= 8'b00110000; // a   **
        1467: q_reg <= 8'b00111100; // b   ****
        1468: q_reg <= 8'b00000000; // c
        1469: q_reg <= 8'b00000000; // d
        1470: q_reg <= 8'b00000000; // e
        1471: q_reg <= 8'b00000000; // f
        // -- code x5c
        1472: q_reg <= 8'b00000000; // 0
        1473: q_reg <= 8'b00000000; // 1
        1474: q_reg <= 8'b00000000; // 2
        1475: q_reg <= 8'b10000000; // 3 *
        1476: q_reg <= 8'b11000000; // 4 **
        1477: q_reg <= 8'b11100000; // 5 ***
        1478: q_reg <= 8'b01110000; // 6  ***
        1479: q_reg <= 8'b00111000; // 7   ***
        1480: q_reg <= 8'b00011100; // 8    ***
        1481: q_reg <= 8'b00001110; // 9     ***
        1482: q_reg <= 8'b00000110; // a      **
        1483: q_reg <= 8'b00000010; // b       *
        1484: q_reg <= 8'b00000000; // c
        1485: q_reg <= 8'b00000000; // d
        1486: q_reg <= 8'b00000000; // e
        1487: q_reg <= 8'b00000000; // f
        // -- code x5d
        1488: q_reg <= 8'b00000000; // 0
        1489: q_reg <= 8'b00000000; // 1
        1490: q_reg <= 8'b00111100; // 2   ****
        1491: q_reg <= 8'b00001100; // 3     **
        1492: q_reg <= 8'b00001100; // 4     **
        1493: q_reg <= 8'b00001100; // 5     **
        1494: q_reg <= 8'b00001100; // 6     **
        1495: q_reg <= 8'b00001100; // 7     **
        1496: q_reg <= 8'b00001100; // 8     **
        1497: q_reg <= 8'b00001100; // 9     **
        1498: q_reg <= 8'b00001100; // a     **
        1499: q_reg <= 8'b00111100; // b   ****
        1500: q_reg <= 8'b00000000; // c
        1501: q_reg <= 8'b00000000; // d
        1502: q_reg <= 8'b00000000; // e
        1503: q_reg <= 8'b00000000; // f
        // -- code x5e
        1504: q_reg <= 8'b00010000; // 0    *
        1505: q_reg <= 8'b00111000; // 1   ***
        1506: q_reg <= 8'b01101100; // 2  ** **
        1507: q_reg <= 8'b11000110; // 3 **   **
        1508: q_reg <= 8'b00000000; // 4
        1509: q_reg <= 8'b00000000; // 5
        1510: q_reg <= 8'b00000000; // 6
        1511: q_reg <= 8'b00000000; // 7
        1512: q_reg <= 8'b00000000; // 8
        1513: q_reg <= 8'b00000000; // 9
        1514: q_reg <= 8'b00000000; // a
        1515: q_reg <= 8'b00000000; // b
        1516: q_reg <= 8'b00000000; // c
        1517: q_reg <= 8'b00000000; // d
        1518: q_reg <= 8'b00000000; // e
        1519: q_reg <= 8'b00000000; // f
        // -- code x5f
        1520: q_reg <= 8'b00000000; // 0
        1521: q_reg <= 8'b00000000; // 1
        1522: q_reg <= 8'b00000000; // 2
        1523: q_reg <= 8'b00000000; // 3
        1524: q_reg <= 8'b00000000; // 4
        1525: q_reg <= 8'b00000000; // 5
        1526: q_reg <= 8'b00000000; // 6
        1527: q_reg <= 8'b00000000; // 7
        1528: q_reg <= 8'b00000000; // 8
        1529: q_reg <= 8'b00000000; // 9
        1530: q_reg <= 8'b00000000; // a
        1531: q_reg <= 8'b00000000; // b
        1532: q_reg <= 8'b00000000; // c
        1533: q_reg <= 8'b11111111; // d ********
        1534: q_reg <= 8'b00000000; // e
        1535: q_reg <= 8'b00000000; // f
        // -- code x60
        1536: q_reg <= 8'b00110000; // 0   **
        1537: q_reg <= 8'b00110000; // 1   **
        1538: q_reg <= 8'b00011000; // 2    **
        1539: q_reg <= 8'b00000000; // 3
        1540: q_reg <= 8'b00000000; // 4
        1541: q_reg <= 8'b00000000; // 5
        1542: q_reg <= 8'b00000000; // 6
        1543: q_reg <= 8'b00000000; // 7
        1544: q_reg <= 8'b00000000; // 8
        1545: q_reg <= 8'b00000000; // 9
        1546: q_reg <= 8'b00000000; // a
        1547: q_reg <= 8'b00000000; // b
        1548: q_reg <= 8'b00000000; // c
        1549: q_reg <= 8'b00000000; // d
        1550: q_reg <= 8'b00000000; // e
        1551: q_reg <= 8'b00000000; // f
        // -- a: code x61
        1552: q_reg <= 8'b00000000; // 0
        1553: q_reg <= 8'b00000000; // 1
        1554: q_reg <= 8'b00000000; // 2
        1555: q_reg <= 8'b00000000; // 3
        1556: q_reg <= 8'b00000000; // 4
        1557: q_reg <= 8'b01111000; // 5  ****
        1558: q_reg <= 8'b00001100; // 6     **
        1559: q_reg <= 8'b01111100; // 7  *****
        1560: q_reg <= 8'b11001100; // 8 **  **
        1561: q_reg <= 8'b11001100; // 9 **  **
        1562: q_reg <= 8'b11001100; // a **  **
        1563: q_reg <= 8'b01110110; // b  *** **
        1564: q_reg <= 8'b00000000; // c
        1565: q_reg <= 8'b00000000; // d
        1566: q_reg <= 8'b00000000; // e
        1567: q_reg <= 8'b00000000; // f
        // -- b: code x62
        1568: q_reg <= 8'b00000000; // 0
        1569: q_reg <= 8'b00000000; // 1
        1570: q_reg <= 8'b11100000; // 2  ***
        1571: q_reg <= 8'b01100000; // 3   **
        1572: q_reg <= 8'b01100000; // 4   **
        1573: q_reg <= 8'b01111000; // 5   ****
        1574: q_reg <= 8'b01101100; // 6   ** **
        1575: q_reg <= 8'b01100110; // 7   **  **
        1576: q_reg <= 8'b01100110; // 8   **  **
        1577: q_reg <= 8'b01100110; // 9   **  **
        1578: q_reg <= 8'b01100110; // a   **  **
        1579: q_reg <= 8'b01111100; // b   *****
        1580: q_reg <= 8'b00000000; // c
        1581: q_reg <= 8'b00000000; // d
        1582: q_reg <= 8'b00000000; // e
        1583: q_reg <= 8'b00000000; // f
        // -- c: code x63
        1584: q_reg <= 8'b00000000; // 0
        1585: q_reg <= 8'b00000000; // 1
        1586: q_reg <= 8'b00000000; // 2
        1587: q_reg <= 8'b00000000; // 3
        1588: q_reg <= 8'b00000000; // 4
        1589: q_reg <= 8'b01111100; // 5  *****
        1590: q_reg <= 8'b11000110; // 6 **   **
        1591: q_reg <= 8'b11000000; // 7 **
        1592: q_reg <= 8'b11000000; // 8 **
        1593: q_reg <= 8'b11000000; // 9 **
        1594: q_reg <= 8'b11000110; // a **   **
        1595: q_reg <= 8'b01111100; // b  *****
        1596: q_reg <= 8'b00000000; // c
        1597: q_reg <= 8'b00000000; // d
        1598: q_reg <= 8'b00000000; // e
        1599: q_reg <= 8'b00000000; // f
        // -- d: code x64
        1600: q_reg <= 8'b00000000; // 0
        1601: q_reg <= 8'b00000000; // 1
        1602: q_reg <= 8'b00011100; // 2    ***
        1603: q_reg <= 8'b00001100; // 3     **
        1604: q_reg <= 8'b00001100; // 4     **
        1605: q_reg <= 8'b00111100; // 5   ****
        1606: q_reg <= 8'b01101100; // 6  ** **
        1607: q_reg <= 8'b11001100; // 7 **  **
        1608: q_reg <= 8'b11001100; // 8 **  **
        1609: q_reg <= 8'b11001100; // 9 **  **
        1610: q_reg <= 8'b11001100; // a **  **
        1611: q_reg <= 8'b01110110; // b  *** **
        1612: q_reg <= 8'b00000000; // c
        1613: q_reg <= 8'b00000000; // d
        1614: q_reg <= 8'b00000000; // e
        1615: q_reg <= 8'b00000000; // f
        // -- e: code x65
        1616: q_reg <= 8'b00000000; // 0
        1617: q_reg <= 8'b00000000; // 1
        1618: q_reg <= 8'b00000000; // 2
        1619: q_reg <= 8'b00000000; // 3
        1620: q_reg <= 8'b00000000; // 4
        1621: q_reg <= 8'b01111100; // 5  *****
        1622: q_reg <= 8'b11000110; // 6 **   **
        1623: q_reg <= 8'b11111110; // 7 *******
        1624: q_reg <= 8'b11000000; // 8 **
        1625: q_reg <= 8'b11000000; // 9 **
        1626: q_reg <= 8'b11000110; // a **   **
        1627: q_reg <= 8'b01111100; // b  *****
        1628: q_reg <= 8'b00000000; // c
        1629: q_reg <= 8'b00000000; // d
        1630: q_reg <= 8'b00000000; // e
        1631: q_reg <= 8'b00000000; // f
        // -- f: code x66
        1632: q_reg <= 8'b00000000; // 0
        1633: q_reg <= 8'b00000000; // 1
        1634: q_reg <= 8'b00111000; // 2   ***
        1635: q_reg <= 8'b01101100; // 3  ** **
        1636: q_reg <= 8'b01100100; // 4  **  *
        1637: q_reg <= 8'b01100000; // 5  **
        1638: q_reg <= 8'b11110000; // 6 ****
        1639: q_reg <= 8'b01100000; // 7  **
        1640: q_reg <= 8'b01100000; // 8  **
        1641: q_reg <= 8'b01100000; // 9  **
        1642: q_reg <= 8'b01100000; // a  **
        1643: q_reg <= 8'b11110000; // b ****
        1644: q_reg <= 8'b00000000; // c
        1645: q_reg <= 8'b00000000; // d
        1646: q_reg <= 8'b00000000; // e
        1647: q_reg <= 8'b00000000; // f
        // -- g: code x67
        1648: q_reg <= 8'b00000000; // 0
        1649: q_reg <= 8'b00000000; // 1
        1650: q_reg <= 8'b00000000; // 2
        1651: q_reg <= 8'b00000000; // 3
        1652: q_reg <= 8'b00000000; // 4
        1653: q_reg <= 8'b01110110; // 5  *** **
        1654: q_reg <= 8'b11001100; // 6 **  **
        1655: q_reg <= 8'b11001100; // 7 **  **
        1656: q_reg <= 8'b11001100; // 8 **  **
        1657: q_reg <= 8'b11001100; // 9 **  **
        1658: q_reg <= 8'b11001100; // a **  **
        1659: q_reg <= 8'b01111100; // b  *****
        1660: q_reg <= 8'b00001100; // c     **
        1661: q_reg <= 8'b11001100; // d **  **
        1662: q_reg <= 8'b01111000; // e  ****
        1663: q_reg <= 8'b00000000; // f
        // -- h: code x68
        1664: q_reg <= 8'b00000000; // 0
        1665: q_reg <= 8'b00000000; // 1
        1666: q_reg <= 8'b11100000; // 2 ***
        1667: q_reg <= 8'b01100000; // 3  **
        1668: q_reg <= 8'b01100000; // 4  **
        1669: q_reg <= 8'b01101100; // 5  ** **
        1670: q_reg <= 8'b01110110; // 6  *** **
        1671: q_reg <= 8'b01100110; // 7  **  **
        1672: q_reg <= 8'b01100110; // 8  **  **
        1673: q_reg <= 8'b01100110; // 9  **  **
        1674: q_reg <= 8'b01100110; // a  **  **
        1675: q_reg <= 8'b11100110; // b ***  **
        1676: q_reg <= 8'b00000000; // c
        1677: q_reg <= 8'b00000000; // d
        1678: q_reg <= 8'b00000000; // e
        1679: q_reg <= 8'b00000000; // f
        // -- i: code x69
        1680: q_reg <= 8'b00000000; // 0
        1681: q_reg <= 8'b00000000; // 1
        1682: q_reg <= 8'b00011000; // 2    **
        1683: q_reg <= 8'b00011000; // 3    **
        1684: q_reg <= 8'b00000000; // 4
        1685: q_reg <= 8'b00111000; // 5   ***
        1686: q_reg <= 8'b00011000; // 6    **
        1687: q_reg <= 8'b00011000; // 7    **
        1688: q_reg <= 8'b00011000; // 8    **
        1689: q_reg <= 8'b00011000; // 9    **
        1690: q_reg <= 8'b00011000; // a    **
        1691: q_reg <= 8'b00111100; // b   ****
        1692: q_reg <= 8'b00000000; // c
        1693: q_reg <= 8'b00000000; // d
        1694: q_reg <= 8'b00000000; // e
        1695: q_reg <= 8'b00000000; // f
        // -- j: code x6a
        1696: q_reg <= 8'b00000000; // 0
        1697: q_reg <= 8'b00000000; // 1
        1698: q_reg <= 8'b00000110; // 2      **
        1699: q_reg <= 8'b00000110; // 3      **
        1700: q_reg <= 8'b00000000; // 4
        1701: q_reg <= 8'b00001110; // 5     ***
        1702: q_reg <= 8'b00000110; // 6      **
        1703: q_reg <= 8'b00000110; // 7      **
        1704: q_reg <= 8'b00000110; // 8      **
        1705: q_reg <= 8'b00000110; // 9      **
        1706: q_reg <= 8'b00000110; // a      **
        1707: q_reg <= 8'b00000110; // b      **
        1708: q_reg <= 8'b01100110; // c  **  **
        1709: q_reg <= 8'b01100110; // d  **  **
        1710: q_reg <= 8'b00111100; // e   ****
        1711: q_reg <= 8'b00000000; // f
        // -- k: code x6b
        1712: q_reg <= 8'b00000000; // 0
        1713: q_reg <= 8'b00000000; // 1
        1714: q_reg <= 8'b11100000; // 2 ***
        1715: q_reg <= 8'b01100000; // 3  **
        1716: q_reg <= 8'b01100000; // 4  **
        1717: q_reg <= 8'b01100110; // 5  **  **
        1718: q_reg <= 8'b01101100; // 6  ** **
        1719: q_reg <= 8'b01111000; // 7  ****
        1720: q_reg <= 8'b01111000; // 8  ****
        1721: q_reg <= 8'b01101100; // 9  ** **
        1722: q_reg <= 8'b01100110; // a  **  **
        1723: q_reg <= 8'b11100110; // b ***  **
        1724: q_reg <= 8'b00000000; // c
        1725: q_reg <= 8'b00000000; // d
        1726: q_reg <= 8'b00000000; // e
        1727: q_reg <= 8'b00000000; // f
        // -- l: code x6c
        1728: q_reg <= 8'b00000000; // 0
        1729: q_reg <= 8'b00000000; // 1
        1730: q_reg <= 8'b00111000; // 2   ***
        1731: q_reg <= 8'b00011000; // 3    **
        1732: q_reg <= 8'b00011000; // 4    **
        1733: q_reg <= 8'b00011000; // 5    **
        1734: q_reg <= 8'b00011000; // 6    **
        1735: q_reg <= 8'b00011000; // 7    **
        1736: q_reg <= 8'b00011000; // 8    **
        1737: q_reg <= 8'b00011000; // 9    **
        1738: q_reg <= 8'b00011000; // a    **
        1739: q_reg <= 8'b00111100; // b   ****
        1740: q_reg <= 8'b00000000; // c
        1741: q_reg <= 8'b00000000; // d
        1742: q_reg <= 8'b00000000; // e
        1743: q_reg <= 8'b00000000; // f
        // -- m: code x6d
        1744: q_reg <= 8'b00000000; // 0
        1745: q_reg <= 8'b00000000; // 1
        1746: q_reg <= 8'b00000000; // 2
        1747: q_reg <= 8'b00000000; // 3
        1748: q_reg <= 8'b00000000; // 4
        1749: q_reg <= 8'b11100110; // 5 ***  **
        1750: q_reg <= 8'b11111111; // 6 ********
        1751: q_reg <= 8'b11011011; // 7 ** ** **
        1752: q_reg <= 8'b11011011; // 8 ** ** **
        1753: q_reg <= 8'b11011011; // 9 ** ** **
        1754: q_reg <= 8'b11011011; // a ** ** **
        1755: q_reg <= 8'b11011011; // b ** ** **
        1756: q_reg <= 8'b00000000; // c
        1757: q_reg <= 8'b00000000; // d
        1758: q_reg <= 8'b00000000; // e
        1759: q_reg <= 8'b00000000; // f
        // -- n: code x6e
        1760: q_reg <= 8'b00000000; // 0
        1761: q_reg <= 8'b00000000; // 1
        1762: q_reg <= 8'b00000000; // 2
        1763: q_reg <= 8'b00000000; // 3
        1764: q_reg <= 8'b00000000; // 4
        1765: q_reg <= 8'b11011100; // 5 ** ***
        1766: q_reg <= 8'b01100110; // 6  **  **
        1767: q_reg <= 8'b01100110; // 7  **  **
        1768: q_reg <= 8'b01100110; // 8  **  **
        1769: q_reg <= 8'b01100110; // 9  **  **
        1770: q_reg <= 8'b01100110; // a  **  **
        1771: q_reg <= 8'b01100110; // b  **  **
        1772: q_reg <= 8'b00000000; // c
        1773: q_reg <= 8'b00000000; // d
        1774: q_reg <= 8'b00000000; // e
        1775: q_reg <= 8'b00000000; // f
        // -- o: code x6f
        1776: q_reg <= 8'b00000000; // 0
        1777: q_reg <= 8'b00000000; // 1
        1778: q_reg <= 8'b00000000; // 2
        1779: q_reg <= 8'b00000000; // 3
        1780: q_reg <= 8'b00000000; // 4
        1781: q_reg <= 8'b01111100; // 5  *****
        1782: q_reg <= 8'b11000110; // 6 **   **
        1783: q_reg <= 8'b11000110; // 7 **   **
        1784: q_reg <= 8'b11000110; // 8 **   **
        1785: q_reg <= 8'b11000110; // 9 **   **
        1786: q_reg <= 8'b11000110; // a **   **
        1787: q_reg <= 8'b01111100; // b  *****
        1788: q_reg <= 8'b00000000; // c
        1789: q_reg <= 8'b00000000; // d
        1790: q_reg <= 8'b00000000; // e
        1791: q_reg <= 8'b00000000; // f
        // -- code x70
        1792: q_reg <= 8'b00000000; // 0
        1793: q_reg <= 8'b00000000; // 1
        1794: q_reg <= 8'b00000000; // 2
        1795: q_reg <= 8'b00000000; // 3
        1796: q_reg <= 8'b00000000; // 4
        1797: q_reg <= 8'b11011100; // 5 ** ***
        1798: q_reg <= 8'b01100110; // 6  **  **
        1799: q_reg <= 8'b01100110; // 7  **  **
        1800: q_reg <= 8'b01100110; // 8  **  **
        1801: q_reg <= 8'b01100110; // 9  **  **
        1802: q_reg <= 8'b01100110; // a  **  **
        1803: q_reg <= 8'b01111100; // b  *****
        1804: q_reg <= 8'b01100000; // c  **
        1805: q_reg <= 8'b01100000; // d  **
        1806: q_reg <= 8'b11110000; // e ****
        1807: q_reg <= 8'b00000000; // f
        // -- code x71
        1808: q_reg <= 8'b00000000; // 0
        1809: q_reg <= 8'b00000000; // 1
        1810: q_reg <= 8'b00000000; // 2
        1811: q_reg <= 8'b00000000; // 3
        1812: q_reg <= 8'b00000000; // 4
        1813: q_reg <= 8'b01110110; // 5  *** **
        1814: q_reg <= 8'b11001100; // 6 **  **
        1815: q_reg <= 8'b11001100; // 7 **  **
        1816: q_reg <= 8'b11001100; // 8 **  **
        1817: q_reg <= 8'b11001100; // 9 **  **
        1818: q_reg <= 8'b11001100; // a **  **
        1819: q_reg <= 8'b01111100; // b  *****
        1820: q_reg <= 8'b00001100; // c     **
        1821: q_reg <= 8'b00001100; // d     **
        1822: q_reg <= 8'b00011110; // e    ****
        1823: q_reg <= 8'b00000000; // f
        // -- code x72
        1824: q_reg <= 8'b00000000; // 0
        1825: q_reg <= 8'b00000000; // 1
        1826: q_reg <= 8'b00000000; // 2
        1827: q_reg <= 8'b00000000; // 3
        1828: q_reg <= 8'b00000000; // 4
        1829: q_reg <= 8'b11011100; // 5 ** ***
        1830: q_reg <= 8'b01110110; // 6  *** **
        1831: q_reg <= 8'b01100110; // 7  **  **
        1832: q_reg <= 8'b01100000; // 8  **
        1833: q_reg <= 8'b01100000; // 9  **
        1834: q_reg <= 8'b01100000; // a  **
        1835: q_reg <= 8'b11110000; // b ****
        1836: q_reg <= 8'b00000000; // c
        1837: q_reg <= 8'b00000000; // d
        1838: q_reg <= 8'b00000000; // e
        1839: q_reg <= 8'b00000000; // f
        // -- code x73
        1840: q_reg <= 8'b00000000; // 0
        1841: q_reg <= 8'b00000000; // 1
        1842: q_reg <= 8'b00000000; // 2
        1843: q_reg <= 8'b00000000; // 3
        1844: q_reg <= 8'b00000000; // 4
        1845: q_reg <= 8'b01111100; // 5  *****
        1846: q_reg <= 8'b11000110; // 6 **   **
        1847: q_reg <= 8'b01100000; // 7  **
        1848: q_reg <= 8'b00111000; // 8   ***
        1849: q_reg <= 8'b00001100; // 9     **
        1850: q_reg <= 8'b11000110; // a **   **
        1851: q_reg <= 8'b01111100; // b  *****
        1852: q_reg <= 8'b00000000; // c
        1853: q_reg <= 8'b00000000; // d
        1854: q_reg <= 8'b00000000; // e
        1855: q_reg <= 8'b00000000; // f
        // -- code x74
        1856: q_reg <= 8'b00000000; // 0
        1857: q_reg <= 8'b00000000; // 1
        1858: q_reg <= 8'b00010000; // 2    *
        1859: q_reg <= 8'b00110000; // 3   **
        1860: q_reg <= 8'b00110000; // 4   **
        1861: q_reg <= 8'b11111100; // 5 ******
        1862: q_reg <= 8'b00110000; // 6   **
        1863: q_reg <= 8'b00110000; // 7   **
        1864: q_reg <= 8'b00110000; // 8   **
        1865: q_reg <= 8'b00110000; // 9   **
        1866: q_reg <= 8'b00110110; // a   ** **
        1867: q_reg <= 8'b00011100; // b    ***
        1868: q_reg <= 8'b00000000; // c
        1869: q_reg <= 8'b00000000; // d
        1870: q_reg <= 8'b00000000; // e
        1871: q_reg <= 8'b00000000; // f
        // -- code x75
        1872: q_reg <= 8'b00000000; // 0
        1873: q_reg <= 8'b00000000; // 1
        1874: q_reg <= 8'b00000000; // 2
        1875: q_reg <= 8'b00000000; // 3
        1876: q_reg <= 8'b00000000; // 4
        1877: q_reg <= 8'b11001100; // 5 **  **
        1878: q_reg <= 8'b11001100; // 6 **  **
        1879: q_reg <= 8'b11001100; // 7 **  **
        1880: q_reg <= 8'b11001100; // 8 **  **
        1881: q_reg <= 8'b11001100; // 9 **  **
        1882: q_reg <= 8'b11001100; // a **  **
        1883: q_reg <= 8'b01110110; // b  *** **
        1884: q_reg <= 8'b00000000; // c
        1885: q_reg <= 8'b00000000; // d
        1886: q_reg <= 8'b00000000; // e
        1887: q_reg <= 8'b00000000; // f
        // -- code x76
        1888: q_reg <= 8'b00000000; // 0
        1889: q_reg <= 8'b00000000; // 1
        1890: q_reg <= 8'b00000000; // 2
        1891: q_reg <= 8'b00000000; // 3
        1892: q_reg <= 8'b00000000; // 4
        1893: q_reg <= 8'b11000011; // 5 **    **
        1894: q_reg <= 8'b11000011; // 6 **    **
        1895: q_reg <= 8'b11000011; // 7 **    **
        1896: q_reg <= 8'b11000011; // 8 **    **
        1897: q_reg <= 8'b01100110; // 9  **  **
        1898: q_reg <= 8'b00111100; // a   ****
        1899: q_reg <= 8'b00011000; // b    **
        1900: q_reg <= 8'b00000000; // c
        1901: q_reg <= 8'b00000000; // d
        1902: q_reg <= 8'b00000000; // e
        1903: q_reg <= 8'b00000000; // f
        // -- code x77
        1904: q_reg <= 8'b00000000; // 0
        1905: q_reg <= 8'b00000000; // 1
        1906: q_reg <= 8'b00000000; // 2
        1907: q_reg <= 8'b00000000; // 3
        1908: q_reg <= 8'b00000000; // 4
        1909: q_reg <= 8'b11000011; // 5 **    **
        1910: q_reg <= 8'b11000011; // 6 **    **
        1911: q_reg <= 8'b11000011; // 7 **    **
        1912: q_reg <= 8'b11011011; // 8 ** ** **
        1913: q_reg <= 8'b11011011; // 9 ** ** **
        1914: q_reg <= 8'b11111111; // a ********
        1915: q_reg <= 8'b01100110; // b  **  **
        1916: q_reg <= 8'b00000000; // c
        1917: q_reg <= 8'b00000000; // d
        1918: q_reg <= 8'b00000000; // e
        1919: q_reg <= 8'b00000000; // f
        // -- code x78
        1920: q_reg <= 8'b00000000; // 0
        1921: q_reg <= 8'b00000000; // 1
        1922: q_reg <= 8'b00000000; // 2
        1923: q_reg <= 8'b00000000; // 3
        1924: q_reg <= 8'b00000000; // 4
        1925: q_reg <= 8'b11000011; // 5 **    **
        1926: q_reg <= 8'b01100110; // 6  **  **
        1927: q_reg <= 8'b00111100; // 7   ****
        1928: q_reg <= 8'b00011000; // 8    **
        1929: q_reg <= 8'b00111100; // 9   ****
        1930: q_reg <= 8'b01100110; // a  **  **
        1931: q_reg <= 8'b11000011; // b **    **
        1932: q_reg <= 8'b00000000; // c
        1933: q_reg <= 8'b00000000; // d
        1934: q_reg <= 8'b00000000; // e
        1935: q_reg <= 8'b00000000; // f
        // -- code x79
        1936: q_reg <= 8'b00000000; // 0
        1937: q_reg <= 8'b00000000; // 1
        1938: q_reg <= 8'b00000000; // 2
        1939: q_reg <= 8'b00000000; // 3
        1940: q_reg <= 8'b00000000; // 4
        1941: q_reg <= 8'b11000110; // 5 **   **
        1942: q_reg <= 8'b11000110; // 6 **   **
        1943: q_reg <= 8'b11000110; // 7 **   **
        1944: q_reg <= 8'b11000110; // 8 **   **
        1945: q_reg <= 8'b11000110; // 9 **   **
        1946: q_reg <= 8'b11000110; // a **   **
        1947: q_reg <= 8'b01111110; // b  ******
        1948: q_reg <= 8'b00000110; // c      **
        1949: q_reg <= 8'b00001100; // d     **
        1950: q_reg <= 8'b11111000; // e *****
        1951: q_reg <= 8'b00000000; // f
        // -- code x7a
        1952: q_reg <= 8'b00000000; // 0
        1953: q_reg <= 8'b00000000; // 1
        1954: q_reg <= 8'b00000000; // 2
        1955: q_reg <= 8'b00000000; // 3
        1956: q_reg <= 8'b00000000; // 4
        1957: q_reg <= 8'b11111110; // 5 *******
        1958: q_reg <= 8'b11001100; // 6 **  **
        1959: q_reg <= 8'b00011000; // 7    **
        1960: q_reg <= 8'b00110000; // 8   **
        1961: q_reg <= 8'b01100000; // 9  **
        1962: q_reg <= 8'b11000110; // a **   **
        1963: q_reg <= 8'b11111110; // b *******
        1964: q_reg <= 8'b00000000; // c
        1965: q_reg <= 8'b00000000; // d
        1966: q_reg <= 8'b00000000; // e
        1967: q_reg <= 8'b00000000; // f
        // -- code x7b
        1968: q_reg <= 8'b00000000; // 0
        1969: q_reg <= 8'b00000000; // 1
        1970: q_reg <= 8'b00001110; // 2     ***
        1971: q_reg <= 8'b00011000; // 3    **
        1972: q_reg <= 8'b00011000; // 4    **
        1973: q_reg <= 8'b00011000; // 5    **
        1974: q_reg <= 8'b01110000; // 6  ***
        1975: q_reg <= 8'b00011000; // 7    **
        1976: q_reg <= 8'b00011000; // 8    **
        1977: q_reg <= 8'b00011000; // 9    **
        1978: q_reg <= 8'b00011000; // a    **
        1979: q_reg <= 8'b00001110; // b     ***
        1980: q_reg <= 8'b00000000; // c
        1981: q_reg <= 8'b00000000; // d
        1982: q_reg <= 8'b00000000; // e
        1983: q_reg <= 8'b00000000; // f
        // -- code x7c
        1984: q_reg <= 8'b00000000; // 0
        1985: q_reg <= 8'b00000000; // 1
        1986: q_reg <= 8'b00011000; // 2    **
        1987: q_reg <= 8'b00011000; // 3    **
        1988: q_reg <= 8'b00011000; // 4    **
        1989: q_reg <= 8'b00011000; // 5    **
        1990: q_reg <= 8'b00000000; // 6
        1991: q_reg <= 8'b00011000; // 7    **
        1992: q_reg <= 8'b00011000; // 8    **
        1993: q_reg <= 8'b00011000; // 9    **
        1994: q_reg <= 8'b00011000; // a    **
        1995: q_reg <= 8'b00011000; // b    **
        1996: q_reg <= 8'b00000000; // c
        1997: q_reg <= 8'b00000000; // d
        1998: q_reg <= 8'b00000000; // e
        1999: q_reg <= 8'b00000000; // f
        // -- code x7d
        2000: q_reg <= 8'b00000000; // 0
        2001: q_reg <= 8'b00000000; // 1
        2002: q_reg <= 8'b01110000; // 2  ***
        2003: q_reg <= 8'b00011000; // 3    **
        2004: q_reg <= 8'b00011000; // 4    **
        2005: q_reg <= 8'b00011000; // 5    **
        2006: q_reg <= 8'b00001110; // 6     ***
        2007: q_reg <= 8'b00011000; // 7    **
        2008: q_reg <= 8'b00011000; // 8    **
        2009: q_reg <= 8'b00011000; // 9    **
        2010: q_reg <= 8'b00011000; // a    **
        2011: q_reg <= 8'b01110000; // b  ***
        2012: q_reg <= 8'b00000000; // c
        2013: q_reg <= 8'b00000000; // d
        2014: q_reg <= 8'b00000000; // e
        2015: q_reg <= 8'b00000000; // f
        // -- code x7e
        2016: q_reg <= 8'b00000000; // 0
        2017: q_reg <= 8'b00000000; // 1
        2018: q_reg <= 8'b01110110; // 2  *** **
        2019: q_reg <= 8'b11011100; // 3 ** ***
        2020: q_reg <= 8'b00000000; // 4
        2021: q_reg <= 8'b00000000; // 5
        2022: q_reg <= 8'b00000000; // 6
        2023: q_reg <= 8'b00000000; // 7
        2024: q_reg <= 8'b00000000; // 8
        2025: q_reg <= 8'b00000000; // 9
        2026: q_reg <= 8'b00000000; // a
        2027: q_reg <= 8'b00000000; // b
        2028: q_reg <= 8'b00000000; // c
        2029: q_reg <= 8'b00000000; // d
        2030: q_reg <= 8'b00000000; // e
        2031: q_reg <= 8'b00000000; // f
        // -- code x7f
        2032: q_reg <= 8'b00000000; // 0
        2033: q_reg <= 8'b00000000; // 1
        2034: q_reg <= 8'b00000000; // 2
        2035: q_reg <= 8'b00000000; // 3
        2036: q_reg <= 8'b00010000; // 4    *
        2037: q_reg <= 8'b00111000; // 5   ***
        2038: q_reg <= 8'b01101100; // 6  ** **
        2039: q_reg <= 8'b11000110; // 7 **   **
        2040: q_reg <= 8'b11000110; // 8 **   **
        2041: q_reg <= 8'b11000110; // 9 **   **
        2042: q_reg <= 8'b11111110; // a *******
        2043: q_reg <= 8'b00000000; // b
        2044: q_reg <= 8'b00000000; // c
        2045: q_reg <= 8'b00000000; // d
        2046: q_reg <= 8'b00000000; // e
        2047: q_reg <= 8'b00000000; // f
    endcase
    q_reg_2 <= q_reg;
end
endmodule
