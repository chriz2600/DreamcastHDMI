
module osc (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
